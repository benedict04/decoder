magic
tech sky130A
magscale 1 2
timestamp 1698989888
<< checkpaint >>
rect -3932 -1804 43932 41516
<< viali >>
rect 38301 21981 38335 22015
rect 38485 21845 38519 21879
rect 1409 21505 1443 21539
rect 20453 21505 20487 21539
rect 38301 21505 38335 21539
rect 1593 21301 1627 21335
rect 19165 21301 19199 21335
rect 38485 21301 38519 21335
rect 19809 20961 19843 20995
rect 1593 20893 1627 20927
rect 19993 20893 20027 20927
rect 38301 20893 38335 20927
rect 19533 20825 19567 20859
rect 20269 20825 20303 20859
rect 1409 20757 1443 20791
rect 19901 20757 19935 20791
rect 38485 20757 38519 20791
rect 19257 20553 19291 20587
rect 20085 20553 20119 20587
rect 20913 20553 20947 20587
rect 19441 20417 19475 20451
rect 20177 20417 20211 20451
rect 20269 20417 20303 20451
rect 20453 20417 20487 20451
rect 20729 20417 20763 20451
rect 19533 20349 19567 20383
rect 19717 20349 19751 20383
rect 20637 20213 20671 20247
rect 38485 20009 38519 20043
rect 1593 19941 1627 19975
rect 22293 19941 22327 19975
rect 18337 19873 18371 19907
rect 18705 19873 18739 19907
rect 1409 19805 1443 19839
rect 18797 19805 18831 19839
rect 19073 19805 19107 19839
rect 21833 19805 21867 19839
rect 22109 19805 22143 19839
rect 38301 19805 38335 19839
rect 21741 19737 21775 19771
rect 18613 19669 18647 19703
rect 20453 19669 20487 19703
rect 22017 19669 22051 19703
rect 18981 19465 19015 19499
rect 19257 19465 19291 19499
rect 21005 19397 21039 19431
rect 1593 19329 1627 19363
rect 18797 19329 18831 19363
rect 19073 19329 19107 19363
rect 19625 19329 19659 19363
rect 19717 19329 19751 19363
rect 19901 19329 19935 19363
rect 20177 19329 20211 19363
rect 20637 19329 20671 19363
rect 21097 19329 21131 19363
rect 21189 19329 21223 19363
rect 38301 19329 38335 19363
rect 20453 19261 20487 19295
rect 19349 19193 19383 19227
rect 1409 19125 1443 19159
rect 38485 19125 38519 19159
rect 21005 18921 21039 18955
rect 1593 18853 1627 18887
rect 19717 18785 19751 18819
rect 1409 18717 1443 18751
rect 19533 18717 19567 18751
rect 20085 18717 20119 18751
rect 21465 18717 21499 18751
rect 38301 18717 38335 18751
rect 20269 18649 20303 18683
rect 20453 18649 20487 18683
rect 20729 18649 20763 18683
rect 20177 18581 20211 18615
rect 20637 18581 20671 18615
rect 20821 18581 20855 18615
rect 22753 18581 22787 18615
rect 38485 18581 38519 18615
rect 19901 18377 19935 18411
rect 20177 18377 20211 18411
rect 19533 18309 19567 18343
rect 19993 18309 20027 18343
rect 19809 18241 19843 18275
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 1950 37562
rect 2002 37510 2014 37562
rect 2066 37510 2078 37562
rect 2130 37510 2142 37562
rect 2194 37510 2206 37562
rect 2258 37510 6950 37562
rect 7002 37510 7014 37562
rect 7066 37510 7078 37562
rect 7130 37510 7142 37562
rect 7194 37510 7206 37562
rect 7258 37510 11950 37562
rect 12002 37510 12014 37562
rect 12066 37510 12078 37562
rect 12130 37510 12142 37562
rect 12194 37510 12206 37562
rect 12258 37510 16950 37562
rect 17002 37510 17014 37562
rect 17066 37510 17078 37562
rect 17130 37510 17142 37562
rect 17194 37510 17206 37562
rect 17258 37510 21950 37562
rect 22002 37510 22014 37562
rect 22066 37510 22078 37562
rect 22130 37510 22142 37562
rect 22194 37510 22206 37562
rect 22258 37510 26950 37562
rect 27002 37510 27014 37562
rect 27066 37510 27078 37562
rect 27130 37510 27142 37562
rect 27194 37510 27206 37562
rect 27258 37510 31950 37562
rect 32002 37510 32014 37562
rect 32066 37510 32078 37562
rect 32130 37510 32142 37562
rect 32194 37510 32206 37562
rect 32258 37510 36950 37562
rect 37002 37510 37014 37562
rect 37066 37510 37078 37562
rect 37130 37510 37142 37562
rect 37194 37510 37206 37562
rect 37258 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 2610 37018
rect 2662 36966 2674 37018
rect 2726 36966 2738 37018
rect 2790 36966 2802 37018
rect 2854 36966 2866 37018
rect 2918 36966 7610 37018
rect 7662 36966 7674 37018
rect 7726 36966 7738 37018
rect 7790 36966 7802 37018
rect 7854 36966 7866 37018
rect 7918 36966 12610 37018
rect 12662 36966 12674 37018
rect 12726 36966 12738 37018
rect 12790 36966 12802 37018
rect 12854 36966 12866 37018
rect 12918 36966 17610 37018
rect 17662 36966 17674 37018
rect 17726 36966 17738 37018
rect 17790 36966 17802 37018
rect 17854 36966 17866 37018
rect 17918 36966 22610 37018
rect 22662 36966 22674 37018
rect 22726 36966 22738 37018
rect 22790 36966 22802 37018
rect 22854 36966 22866 37018
rect 22918 36966 27610 37018
rect 27662 36966 27674 37018
rect 27726 36966 27738 37018
rect 27790 36966 27802 37018
rect 27854 36966 27866 37018
rect 27918 36966 32610 37018
rect 32662 36966 32674 37018
rect 32726 36966 32738 37018
rect 32790 36966 32802 37018
rect 32854 36966 32866 37018
rect 32918 36966 37610 37018
rect 37662 36966 37674 37018
rect 37726 36966 37738 37018
rect 37790 36966 37802 37018
rect 37854 36966 37866 37018
rect 37918 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 1950 36474
rect 2002 36422 2014 36474
rect 2066 36422 2078 36474
rect 2130 36422 2142 36474
rect 2194 36422 2206 36474
rect 2258 36422 6950 36474
rect 7002 36422 7014 36474
rect 7066 36422 7078 36474
rect 7130 36422 7142 36474
rect 7194 36422 7206 36474
rect 7258 36422 11950 36474
rect 12002 36422 12014 36474
rect 12066 36422 12078 36474
rect 12130 36422 12142 36474
rect 12194 36422 12206 36474
rect 12258 36422 16950 36474
rect 17002 36422 17014 36474
rect 17066 36422 17078 36474
rect 17130 36422 17142 36474
rect 17194 36422 17206 36474
rect 17258 36422 21950 36474
rect 22002 36422 22014 36474
rect 22066 36422 22078 36474
rect 22130 36422 22142 36474
rect 22194 36422 22206 36474
rect 22258 36422 26950 36474
rect 27002 36422 27014 36474
rect 27066 36422 27078 36474
rect 27130 36422 27142 36474
rect 27194 36422 27206 36474
rect 27258 36422 31950 36474
rect 32002 36422 32014 36474
rect 32066 36422 32078 36474
rect 32130 36422 32142 36474
rect 32194 36422 32206 36474
rect 32258 36422 36950 36474
rect 37002 36422 37014 36474
rect 37066 36422 37078 36474
rect 37130 36422 37142 36474
rect 37194 36422 37206 36474
rect 37258 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 2610 35930
rect 2662 35878 2674 35930
rect 2726 35878 2738 35930
rect 2790 35878 2802 35930
rect 2854 35878 2866 35930
rect 2918 35878 7610 35930
rect 7662 35878 7674 35930
rect 7726 35878 7738 35930
rect 7790 35878 7802 35930
rect 7854 35878 7866 35930
rect 7918 35878 12610 35930
rect 12662 35878 12674 35930
rect 12726 35878 12738 35930
rect 12790 35878 12802 35930
rect 12854 35878 12866 35930
rect 12918 35878 17610 35930
rect 17662 35878 17674 35930
rect 17726 35878 17738 35930
rect 17790 35878 17802 35930
rect 17854 35878 17866 35930
rect 17918 35878 22610 35930
rect 22662 35878 22674 35930
rect 22726 35878 22738 35930
rect 22790 35878 22802 35930
rect 22854 35878 22866 35930
rect 22918 35878 27610 35930
rect 27662 35878 27674 35930
rect 27726 35878 27738 35930
rect 27790 35878 27802 35930
rect 27854 35878 27866 35930
rect 27918 35878 32610 35930
rect 32662 35878 32674 35930
rect 32726 35878 32738 35930
rect 32790 35878 32802 35930
rect 32854 35878 32866 35930
rect 32918 35878 37610 35930
rect 37662 35878 37674 35930
rect 37726 35878 37738 35930
rect 37790 35878 37802 35930
rect 37854 35878 37866 35930
rect 37918 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 1950 35386
rect 2002 35334 2014 35386
rect 2066 35334 2078 35386
rect 2130 35334 2142 35386
rect 2194 35334 2206 35386
rect 2258 35334 6950 35386
rect 7002 35334 7014 35386
rect 7066 35334 7078 35386
rect 7130 35334 7142 35386
rect 7194 35334 7206 35386
rect 7258 35334 11950 35386
rect 12002 35334 12014 35386
rect 12066 35334 12078 35386
rect 12130 35334 12142 35386
rect 12194 35334 12206 35386
rect 12258 35334 16950 35386
rect 17002 35334 17014 35386
rect 17066 35334 17078 35386
rect 17130 35334 17142 35386
rect 17194 35334 17206 35386
rect 17258 35334 21950 35386
rect 22002 35334 22014 35386
rect 22066 35334 22078 35386
rect 22130 35334 22142 35386
rect 22194 35334 22206 35386
rect 22258 35334 26950 35386
rect 27002 35334 27014 35386
rect 27066 35334 27078 35386
rect 27130 35334 27142 35386
rect 27194 35334 27206 35386
rect 27258 35334 31950 35386
rect 32002 35334 32014 35386
rect 32066 35334 32078 35386
rect 32130 35334 32142 35386
rect 32194 35334 32206 35386
rect 32258 35334 36950 35386
rect 37002 35334 37014 35386
rect 37066 35334 37078 35386
rect 37130 35334 37142 35386
rect 37194 35334 37206 35386
rect 37258 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 2610 34842
rect 2662 34790 2674 34842
rect 2726 34790 2738 34842
rect 2790 34790 2802 34842
rect 2854 34790 2866 34842
rect 2918 34790 7610 34842
rect 7662 34790 7674 34842
rect 7726 34790 7738 34842
rect 7790 34790 7802 34842
rect 7854 34790 7866 34842
rect 7918 34790 12610 34842
rect 12662 34790 12674 34842
rect 12726 34790 12738 34842
rect 12790 34790 12802 34842
rect 12854 34790 12866 34842
rect 12918 34790 17610 34842
rect 17662 34790 17674 34842
rect 17726 34790 17738 34842
rect 17790 34790 17802 34842
rect 17854 34790 17866 34842
rect 17918 34790 22610 34842
rect 22662 34790 22674 34842
rect 22726 34790 22738 34842
rect 22790 34790 22802 34842
rect 22854 34790 22866 34842
rect 22918 34790 27610 34842
rect 27662 34790 27674 34842
rect 27726 34790 27738 34842
rect 27790 34790 27802 34842
rect 27854 34790 27866 34842
rect 27918 34790 32610 34842
rect 32662 34790 32674 34842
rect 32726 34790 32738 34842
rect 32790 34790 32802 34842
rect 32854 34790 32866 34842
rect 32918 34790 37610 34842
rect 37662 34790 37674 34842
rect 37726 34790 37738 34842
rect 37790 34790 37802 34842
rect 37854 34790 37866 34842
rect 37918 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 1950 34298
rect 2002 34246 2014 34298
rect 2066 34246 2078 34298
rect 2130 34246 2142 34298
rect 2194 34246 2206 34298
rect 2258 34246 6950 34298
rect 7002 34246 7014 34298
rect 7066 34246 7078 34298
rect 7130 34246 7142 34298
rect 7194 34246 7206 34298
rect 7258 34246 11950 34298
rect 12002 34246 12014 34298
rect 12066 34246 12078 34298
rect 12130 34246 12142 34298
rect 12194 34246 12206 34298
rect 12258 34246 16950 34298
rect 17002 34246 17014 34298
rect 17066 34246 17078 34298
rect 17130 34246 17142 34298
rect 17194 34246 17206 34298
rect 17258 34246 21950 34298
rect 22002 34246 22014 34298
rect 22066 34246 22078 34298
rect 22130 34246 22142 34298
rect 22194 34246 22206 34298
rect 22258 34246 26950 34298
rect 27002 34246 27014 34298
rect 27066 34246 27078 34298
rect 27130 34246 27142 34298
rect 27194 34246 27206 34298
rect 27258 34246 31950 34298
rect 32002 34246 32014 34298
rect 32066 34246 32078 34298
rect 32130 34246 32142 34298
rect 32194 34246 32206 34298
rect 32258 34246 36950 34298
rect 37002 34246 37014 34298
rect 37066 34246 37078 34298
rect 37130 34246 37142 34298
rect 37194 34246 37206 34298
rect 37258 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 2610 33754
rect 2662 33702 2674 33754
rect 2726 33702 2738 33754
rect 2790 33702 2802 33754
rect 2854 33702 2866 33754
rect 2918 33702 7610 33754
rect 7662 33702 7674 33754
rect 7726 33702 7738 33754
rect 7790 33702 7802 33754
rect 7854 33702 7866 33754
rect 7918 33702 12610 33754
rect 12662 33702 12674 33754
rect 12726 33702 12738 33754
rect 12790 33702 12802 33754
rect 12854 33702 12866 33754
rect 12918 33702 17610 33754
rect 17662 33702 17674 33754
rect 17726 33702 17738 33754
rect 17790 33702 17802 33754
rect 17854 33702 17866 33754
rect 17918 33702 22610 33754
rect 22662 33702 22674 33754
rect 22726 33702 22738 33754
rect 22790 33702 22802 33754
rect 22854 33702 22866 33754
rect 22918 33702 27610 33754
rect 27662 33702 27674 33754
rect 27726 33702 27738 33754
rect 27790 33702 27802 33754
rect 27854 33702 27866 33754
rect 27918 33702 32610 33754
rect 32662 33702 32674 33754
rect 32726 33702 32738 33754
rect 32790 33702 32802 33754
rect 32854 33702 32866 33754
rect 32918 33702 37610 33754
rect 37662 33702 37674 33754
rect 37726 33702 37738 33754
rect 37790 33702 37802 33754
rect 37854 33702 37866 33754
rect 37918 33702 38824 33754
rect 1104 33680 38824 33702
rect 1104 33210 38824 33232
rect 1104 33158 1950 33210
rect 2002 33158 2014 33210
rect 2066 33158 2078 33210
rect 2130 33158 2142 33210
rect 2194 33158 2206 33210
rect 2258 33158 6950 33210
rect 7002 33158 7014 33210
rect 7066 33158 7078 33210
rect 7130 33158 7142 33210
rect 7194 33158 7206 33210
rect 7258 33158 11950 33210
rect 12002 33158 12014 33210
rect 12066 33158 12078 33210
rect 12130 33158 12142 33210
rect 12194 33158 12206 33210
rect 12258 33158 16950 33210
rect 17002 33158 17014 33210
rect 17066 33158 17078 33210
rect 17130 33158 17142 33210
rect 17194 33158 17206 33210
rect 17258 33158 21950 33210
rect 22002 33158 22014 33210
rect 22066 33158 22078 33210
rect 22130 33158 22142 33210
rect 22194 33158 22206 33210
rect 22258 33158 26950 33210
rect 27002 33158 27014 33210
rect 27066 33158 27078 33210
rect 27130 33158 27142 33210
rect 27194 33158 27206 33210
rect 27258 33158 31950 33210
rect 32002 33158 32014 33210
rect 32066 33158 32078 33210
rect 32130 33158 32142 33210
rect 32194 33158 32206 33210
rect 32258 33158 36950 33210
rect 37002 33158 37014 33210
rect 37066 33158 37078 33210
rect 37130 33158 37142 33210
rect 37194 33158 37206 33210
rect 37258 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 2610 32666
rect 2662 32614 2674 32666
rect 2726 32614 2738 32666
rect 2790 32614 2802 32666
rect 2854 32614 2866 32666
rect 2918 32614 7610 32666
rect 7662 32614 7674 32666
rect 7726 32614 7738 32666
rect 7790 32614 7802 32666
rect 7854 32614 7866 32666
rect 7918 32614 12610 32666
rect 12662 32614 12674 32666
rect 12726 32614 12738 32666
rect 12790 32614 12802 32666
rect 12854 32614 12866 32666
rect 12918 32614 17610 32666
rect 17662 32614 17674 32666
rect 17726 32614 17738 32666
rect 17790 32614 17802 32666
rect 17854 32614 17866 32666
rect 17918 32614 22610 32666
rect 22662 32614 22674 32666
rect 22726 32614 22738 32666
rect 22790 32614 22802 32666
rect 22854 32614 22866 32666
rect 22918 32614 27610 32666
rect 27662 32614 27674 32666
rect 27726 32614 27738 32666
rect 27790 32614 27802 32666
rect 27854 32614 27866 32666
rect 27918 32614 32610 32666
rect 32662 32614 32674 32666
rect 32726 32614 32738 32666
rect 32790 32614 32802 32666
rect 32854 32614 32866 32666
rect 32918 32614 37610 32666
rect 37662 32614 37674 32666
rect 37726 32614 37738 32666
rect 37790 32614 37802 32666
rect 37854 32614 37866 32666
rect 37918 32614 38824 32666
rect 1104 32592 38824 32614
rect 1104 32122 38824 32144
rect 1104 32070 1950 32122
rect 2002 32070 2014 32122
rect 2066 32070 2078 32122
rect 2130 32070 2142 32122
rect 2194 32070 2206 32122
rect 2258 32070 6950 32122
rect 7002 32070 7014 32122
rect 7066 32070 7078 32122
rect 7130 32070 7142 32122
rect 7194 32070 7206 32122
rect 7258 32070 11950 32122
rect 12002 32070 12014 32122
rect 12066 32070 12078 32122
rect 12130 32070 12142 32122
rect 12194 32070 12206 32122
rect 12258 32070 16950 32122
rect 17002 32070 17014 32122
rect 17066 32070 17078 32122
rect 17130 32070 17142 32122
rect 17194 32070 17206 32122
rect 17258 32070 21950 32122
rect 22002 32070 22014 32122
rect 22066 32070 22078 32122
rect 22130 32070 22142 32122
rect 22194 32070 22206 32122
rect 22258 32070 26950 32122
rect 27002 32070 27014 32122
rect 27066 32070 27078 32122
rect 27130 32070 27142 32122
rect 27194 32070 27206 32122
rect 27258 32070 31950 32122
rect 32002 32070 32014 32122
rect 32066 32070 32078 32122
rect 32130 32070 32142 32122
rect 32194 32070 32206 32122
rect 32258 32070 36950 32122
rect 37002 32070 37014 32122
rect 37066 32070 37078 32122
rect 37130 32070 37142 32122
rect 37194 32070 37206 32122
rect 37258 32070 38824 32122
rect 1104 32048 38824 32070
rect 1104 31578 38824 31600
rect 1104 31526 2610 31578
rect 2662 31526 2674 31578
rect 2726 31526 2738 31578
rect 2790 31526 2802 31578
rect 2854 31526 2866 31578
rect 2918 31526 7610 31578
rect 7662 31526 7674 31578
rect 7726 31526 7738 31578
rect 7790 31526 7802 31578
rect 7854 31526 7866 31578
rect 7918 31526 12610 31578
rect 12662 31526 12674 31578
rect 12726 31526 12738 31578
rect 12790 31526 12802 31578
rect 12854 31526 12866 31578
rect 12918 31526 17610 31578
rect 17662 31526 17674 31578
rect 17726 31526 17738 31578
rect 17790 31526 17802 31578
rect 17854 31526 17866 31578
rect 17918 31526 22610 31578
rect 22662 31526 22674 31578
rect 22726 31526 22738 31578
rect 22790 31526 22802 31578
rect 22854 31526 22866 31578
rect 22918 31526 27610 31578
rect 27662 31526 27674 31578
rect 27726 31526 27738 31578
rect 27790 31526 27802 31578
rect 27854 31526 27866 31578
rect 27918 31526 32610 31578
rect 32662 31526 32674 31578
rect 32726 31526 32738 31578
rect 32790 31526 32802 31578
rect 32854 31526 32866 31578
rect 32918 31526 37610 31578
rect 37662 31526 37674 31578
rect 37726 31526 37738 31578
rect 37790 31526 37802 31578
rect 37854 31526 37866 31578
rect 37918 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 1950 31034
rect 2002 30982 2014 31034
rect 2066 30982 2078 31034
rect 2130 30982 2142 31034
rect 2194 30982 2206 31034
rect 2258 30982 6950 31034
rect 7002 30982 7014 31034
rect 7066 30982 7078 31034
rect 7130 30982 7142 31034
rect 7194 30982 7206 31034
rect 7258 30982 11950 31034
rect 12002 30982 12014 31034
rect 12066 30982 12078 31034
rect 12130 30982 12142 31034
rect 12194 30982 12206 31034
rect 12258 30982 16950 31034
rect 17002 30982 17014 31034
rect 17066 30982 17078 31034
rect 17130 30982 17142 31034
rect 17194 30982 17206 31034
rect 17258 30982 21950 31034
rect 22002 30982 22014 31034
rect 22066 30982 22078 31034
rect 22130 30982 22142 31034
rect 22194 30982 22206 31034
rect 22258 30982 26950 31034
rect 27002 30982 27014 31034
rect 27066 30982 27078 31034
rect 27130 30982 27142 31034
rect 27194 30982 27206 31034
rect 27258 30982 31950 31034
rect 32002 30982 32014 31034
rect 32066 30982 32078 31034
rect 32130 30982 32142 31034
rect 32194 30982 32206 31034
rect 32258 30982 36950 31034
rect 37002 30982 37014 31034
rect 37066 30982 37078 31034
rect 37130 30982 37142 31034
rect 37194 30982 37206 31034
rect 37258 30982 38824 31034
rect 1104 30960 38824 30982
rect 1104 30490 38824 30512
rect 1104 30438 2610 30490
rect 2662 30438 2674 30490
rect 2726 30438 2738 30490
rect 2790 30438 2802 30490
rect 2854 30438 2866 30490
rect 2918 30438 7610 30490
rect 7662 30438 7674 30490
rect 7726 30438 7738 30490
rect 7790 30438 7802 30490
rect 7854 30438 7866 30490
rect 7918 30438 12610 30490
rect 12662 30438 12674 30490
rect 12726 30438 12738 30490
rect 12790 30438 12802 30490
rect 12854 30438 12866 30490
rect 12918 30438 17610 30490
rect 17662 30438 17674 30490
rect 17726 30438 17738 30490
rect 17790 30438 17802 30490
rect 17854 30438 17866 30490
rect 17918 30438 22610 30490
rect 22662 30438 22674 30490
rect 22726 30438 22738 30490
rect 22790 30438 22802 30490
rect 22854 30438 22866 30490
rect 22918 30438 27610 30490
rect 27662 30438 27674 30490
rect 27726 30438 27738 30490
rect 27790 30438 27802 30490
rect 27854 30438 27866 30490
rect 27918 30438 32610 30490
rect 32662 30438 32674 30490
rect 32726 30438 32738 30490
rect 32790 30438 32802 30490
rect 32854 30438 32866 30490
rect 32918 30438 37610 30490
rect 37662 30438 37674 30490
rect 37726 30438 37738 30490
rect 37790 30438 37802 30490
rect 37854 30438 37866 30490
rect 37918 30438 38824 30490
rect 1104 30416 38824 30438
rect 1104 29946 38824 29968
rect 1104 29894 1950 29946
rect 2002 29894 2014 29946
rect 2066 29894 2078 29946
rect 2130 29894 2142 29946
rect 2194 29894 2206 29946
rect 2258 29894 6950 29946
rect 7002 29894 7014 29946
rect 7066 29894 7078 29946
rect 7130 29894 7142 29946
rect 7194 29894 7206 29946
rect 7258 29894 11950 29946
rect 12002 29894 12014 29946
rect 12066 29894 12078 29946
rect 12130 29894 12142 29946
rect 12194 29894 12206 29946
rect 12258 29894 16950 29946
rect 17002 29894 17014 29946
rect 17066 29894 17078 29946
rect 17130 29894 17142 29946
rect 17194 29894 17206 29946
rect 17258 29894 21950 29946
rect 22002 29894 22014 29946
rect 22066 29894 22078 29946
rect 22130 29894 22142 29946
rect 22194 29894 22206 29946
rect 22258 29894 26950 29946
rect 27002 29894 27014 29946
rect 27066 29894 27078 29946
rect 27130 29894 27142 29946
rect 27194 29894 27206 29946
rect 27258 29894 31950 29946
rect 32002 29894 32014 29946
rect 32066 29894 32078 29946
rect 32130 29894 32142 29946
rect 32194 29894 32206 29946
rect 32258 29894 36950 29946
rect 37002 29894 37014 29946
rect 37066 29894 37078 29946
rect 37130 29894 37142 29946
rect 37194 29894 37206 29946
rect 37258 29894 38824 29946
rect 1104 29872 38824 29894
rect 1104 29402 38824 29424
rect 1104 29350 2610 29402
rect 2662 29350 2674 29402
rect 2726 29350 2738 29402
rect 2790 29350 2802 29402
rect 2854 29350 2866 29402
rect 2918 29350 7610 29402
rect 7662 29350 7674 29402
rect 7726 29350 7738 29402
rect 7790 29350 7802 29402
rect 7854 29350 7866 29402
rect 7918 29350 12610 29402
rect 12662 29350 12674 29402
rect 12726 29350 12738 29402
rect 12790 29350 12802 29402
rect 12854 29350 12866 29402
rect 12918 29350 17610 29402
rect 17662 29350 17674 29402
rect 17726 29350 17738 29402
rect 17790 29350 17802 29402
rect 17854 29350 17866 29402
rect 17918 29350 22610 29402
rect 22662 29350 22674 29402
rect 22726 29350 22738 29402
rect 22790 29350 22802 29402
rect 22854 29350 22866 29402
rect 22918 29350 27610 29402
rect 27662 29350 27674 29402
rect 27726 29350 27738 29402
rect 27790 29350 27802 29402
rect 27854 29350 27866 29402
rect 27918 29350 32610 29402
rect 32662 29350 32674 29402
rect 32726 29350 32738 29402
rect 32790 29350 32802 29402
rect 32854 29350 32866 29402
rect 32918 29350 37610 29402
rect 37662 29350 37674 29402
rect 37726 29350 37738 29402
rect 37790 29350 37802 29402
rect 37854 29350 37866 29402
rect 37918 29350 38824 29402
rect 1104 29328 38824 29350
rect 1104 28858 38824 28880
rect 1104 28806 1950 28858
rect 2002 28806 2014 28858
rect 2066 28806 2078 28858
rect 2130 28806 2142 28858
rect 2194 28806 2206 28858
rect 2258 28806 6950 28858
rect 7002 28806 7014 28858
rect 7066 28806 7078 28858
rect 7130 28806 7142 28858
rect 7194 28806 7206 28858
rect 7258 28806 11950 28858
rect 12002 28806 12014 28858
rect 12066 28806 12078 28858
rect 12130 28806 12142 28858
rect 12194 28806 12206 28858
rect 12258 28806 16950 28858
rect 17002 28806 17014 28858
rect 17066 28806 17078 28858
rect 17130 28806 17142 28858
rect 17194 28806 17206 28858
rect 17258 28806 21950 28858
rect 22002 28806 22014 28858
rect 22066 28806 22078 28858
rect 22130 28806 22142 28858
rect 22194 28806 22206 28858
rect 22258 28806 26950 28858
rect 27002 28806 27014 28858
rect 27066 28806 27078 28858
rect 27130 28806 27142 28858
rect 27194 28806 27206 28858
rect 27258 28806 31950 28858
rect 32002 28806 32014 28858
rect 32066 28806 32078 28858
rect 32130 28806 32142 28858
rect 32194 28806 32206 28858
rect 32258 28806 36950 28858
rect 37002 28806 37014 28858
rect 37066 28806 37078 28858
rect 37130 28806 37142 28858
rect 37194 28806 37206 28858
rect 37258 28806 38824 28858
rect 1104 28784 38824 28806
rect 1104 28314 38824 28336
rect 1104 28262 2610 28314
rect 2662 28262 2674 28314
rect 2726 28262 2738 28314
rect 2790 28262 2802 28314
rect 2854 28262 2866 28314
rect 2918 28262 7610 28314
rect 7662 28262 7674 28314
rect 7726 28262 7738 28314
rect 7790 28262 7802 28314
rect 7854 28262 7866 28314
rect 7918 28262 12610 28314
rect 12662 28262 12674 28314
rect 12726 28262 12738 28314
rect 12790 28262 12802 28314
rect 12854 28262 12866 28314
rect 12918 28262 17610 28314
rect 17662 28262 17674 28314
rect 17726 28262 17738 28314
rect 17790 28262 17802 28314
rect 17854 28262 17866 28314
rect 17918 28262 22610 28314
rect 22662 28262 22674 28314
rect 22726 28262 22738 28314
rect 22790 28262 22802 28314
rect 22854 28262 22866 28314
rect 22918 28262 27610 28314
rect 27662 28262 27674 28314
rect 27726 28262 27738 28314
rect 27790 28262 27802 28314
rect 27854 28262 27866 28314
rect 27918 28262 32610 28314
rect 32662 28262 32674 28314
rect 32726 28262 32738 28314
rect 32790 28262 32802 28314
rect 32854 28262 32866 28314
rect 32918 28262 37610 28314
rect 37662 28262 37674 28314
rect 37726 28262 37738 28314
rect 37790 28262 37802 28314
rect 37854 28262 37866 28314
rect 37918 28262 38824 28314
rect 1104 28240 38824 28262
rect 1104 27770 38824 27792
rect 1104 27718 1950 27770
rect 2002 27718 2014 27770
rect 2066 27718 2078 27770
rect 2130 27718 2142 27770
rect 2194 27718 2206 27770
rect 2258 27718 6950 27770
rect 7002 27718 7014 27770
rect 7066 27718 7078 27770
rect 7130 27718 7142 27770
rect 7194 27718 7206 27770
rect 7258 27718 11950 27770
rect 12002 27718 12014 27770
rect 12066 27718 12078 27770
rect 12130 27718 12142 27770
rect 12194 27718 12206 27770
rect 12258 27718 16950 27770
rect 17002 27718 17014 27770
rect 17066 27718 17078 27770
rect 17130 27718 17142 27770
rect 17194 27718 17206 27770
rect 17258 27718 21950 27770
rect 22002 27718 22014 27770
rect 22066 27718 22078 27770
rect 22130 27718 22142 27770
rect 22194 27718 22206 27770
rect 22258 27718 26950 27770
rect 27002 27718 27014 27770
rect 27066 27718 27078 27770
rect 27130 27718 27142 27770
rect 27194 27718 27206 27770
rect 27258 27718 31950 27770
rect 32002 27718 32014 27770
rect 32066 27718 32078 27770
rect 32130 27718 32142 27770
rect 32194 27718 32206 27770
rect 32258 27718 36950 27770
rect 37002 27718 37014 27770
rect 37066 27718 37078 27770
rect 37130 27718 37142 27770
rect 37194 27718 37206 27770
rect 37258 27718 38824 27770
rect 1104 27696 38824 27718
rect 1104 27226 38824 27248
rect 1104 27174 2610 27226
rect 2662 27174 2674 27226
rect 2726 27174 2738 27226
rect 2790 27174 2802 27226
rect 2854 27174 2866 27226
rect 2918 27174 7610 27226
rect 7662 27174 7674 27226
rect 7726 27174 7738 27226
rect 7790 27174 7802 27226
rect 7854 27174 7866 27226
rect 7918 27174 12610 27226
rect 12662 27174 12674 27226
rect 12726 27174 12738 27226
rect 12790 27174 12802 27226
rect 12854 27174 12866 27226
rect 12918 27174 17610 27226
rect 17662 27174 17674 27226
rect 17726 27174 17738 27226
rect 17790 27174 17802 27226
rect 17854 27174 17866 27226
rect 17918 27174 22610 27226
rect 22662 27174 22674 27226
rect 22726 27174 22738 27226
rect 22790 27174 22802 27226
rect 22854 27174 22866 27226
rect 22918 27174 27610 27226
rect 27662 27174 27674 27226
rect 27726 27174 27738 27226
rect 27790 27174 27802 27226
rect 27854 27174 27866 27226
rect 27918 27174 32610 27226
rect 32662 27174 32674 27226
rect 32726 27174 32738 27226
rect 32790 27174 32802 27226
rect 32854 27174 32866 27226
rect 32918 27174 37610 27226
rect 37662 27174 37674 27226
rect 37726 27174 37738 27226
rect 37790 27174 37802 27226
rect 37854 27174 37866 27226
rect 37918 27174 38824 27226
rect 1104 27152 38824 27174
rect 1104 26682 38824 26704
rect 1104 26630 1950 26682
rect 2002 26630 2014 26682
rect 2066 26630 2078 26682
rect 2130 26630 2142 26682
rect 2194 26630 2206 26682
rect 2258 26630 6950 26682
rect 7002 26630 7014 26682
rect 7066 26630 7078 26682
rect 7130 26630 7142 26682
rect 7194 26630 7206 26682
rect 7258 26630 11950 26682
rect 12002 26630 12014 26682
rect 12066 26630 12078 26682
rect 12130 26630 12142 26682
rect 12194 26630 12206 26682
rect 12258 26630 16950 26682
rect 17002 26630 17014 26682
rect 17066 26630 17078 26682
rect 17130 26630 17142 26682
rect 17194 26630 17206 26682
rect 17258 26630 21950 26682
rect 22002 26630 22014 26682
rect 22066 26630 22078 26682
rect 22130 26630 22142 26682
rect 22194 26630 22206 26682
rect 22258 26630 26950 26682
rect 27002 26630 27014 26682
rect 27066 26630 27078 26682
rect 27130 26630 27142 26682
rect 27194 26630 27206 26682
rect 27258 26630 31950 26682
rect 32002 26630 32014 26682
rect 32066 26630 32078 26682
rect 32130 26630 32142 26682
rect 32194 26630 32206 26682
rect 32258 26630 36950 26682
rect 37002 26630 37014 26682
rect 37066 26630 37078 26682
rect 37130 26630 37142 26682
rect 37194 26630 37206 26682
rect 37258 26630 38824 26682
rect 1104 26608 38824 26630
rect 1104 26138 38824 26160
rect 1104 26086 2610 26138
rect 2662 26086 2674 26138
rect 2726 26086 2738 26138
rect 2790 26086 2802 26138
rect 2854 26086 2866 26138
rect 2918 26086 7610 26138
rect 7662 26086 7674 26138
rect 7726 26086 7738 26138
rect 7790 26086 7802 26138
rect 7854 26086 7866 26138
rect 7918 26086 12610 26138
rect 12662 26086 12674 26138
rect 12726 26086 12738 26138
rect 12790 26086 12802 26138
rect 12854 26086 12866 26138
rect 12918 26086 17610 26138
rect 17662 26086 17674 26138
rect 17726 26086 17738 26138
rect 17790 26086 17802 26138
rect 17854 26086 17866 26138
rect 17918 26086 22610 26138
rect 22662 26086 22674 26138
rect 22726 26086 22738 26138
rect 22790 26086 22802 26138
rect 22854 26086 22866 26138
rect 22918 26086 27610 26138
rect 27662 26086 27674 26138
rect 27726 26086 27738 26138
rect 27790 26086 27802 26138
rect 27854 26086 27866 26138
rect 27918 26086 32610 26138
rect 32662 26086 32674 26138
rect 32726 26086 32738 26138
rect 32790 26086 32802 26138
rect 32854 26086 32866 26138
rect 32918 26086 37610 26138
rect 37662 26086 37674 26138
rect 37726 26086 37738 26138
rect 37790 26086 37802 26138
rect 37854 26086 37866 26138
rect 37918 26086 38824 26138
rect 1104 26064 38824 26086
rect 1104 25594 38824 25616
rect 1104 25542 1950 25594
rect 2002 25542 2014 25594
rect 2066 25542 2078 25594
rect 2130 25542 2142 25594
rect 2194 25542 2206 25594
rect 2258 25542 6950 25594
rect 7002 25542 7014 25594
rect 7066 25542 7078 25594
rect 7130 25542 7142 25594
rect 7194 25542 7206 25594
rect 7258 25542 11950 25594
rect 12002 25542 12014 25594
rect 12066 25542 12078 25594
rect 12130 25542 12142 25594
rect 12194 25542 12206 25594
rect 12258 25542 16950 25594
rect 17002 25542 17014 25594
rect 17066 25542 17078 25594
rect 17130 25542 17142 25594
rect 17194 25542 17206 25594
rect 17258 25542 21950 25594
rect 22002 25542 22014 25594
rect 22066 25542 22078 25594
rect 22130 25542 22142 25594
rect 22194 25542 22206 25594
rect 22258 25542 26950 25594
rect 27002 25542 27014 25594
rect 27066 25542 27078 25594
rect 27130 25542 27142 25594
rect 27194 25542 27206 25594
rect 27258 25542 31950 25594
rect 32002 25542 32014 25594
rect 32066 25542 32078 25594
rect 32130 25542 32142 25594
rect 32194 25542 32206 25594
rect 32258 25542 36950 25594
rect 37002 25542 37014 25594
rect 37066 25542 37078 25594
rect 37130 25542 37142 25594
rect 37194 25542 37206 25594
rect 37258 25542 38824 25594
rect 1104 25520 38824 25542
rect 1104 25050 38824 25072
rect 1104 24998 2610 25050
rect 2662 24998 2674 25050
rect 2726 24998 2738 25050
rect 2790 24998 2802 25050
rect 2854 24998 2866 25050
rect 2918 24998 7610 25050
rect 7662 24998 7674 25050
rect 7726 24998 7738 25050
rect 7790 24998 7802 25050
rect 7854 24998 7866 25050
rect 7918 24998 12610 25050
rect 12662 24998 12674 25050
rect 12726 24998 12738 25050
rect 12790 24998 12802 25050
rect 12854 24998 12866 25050
rect 12918 24998 17610 25050
rect 17662 24998 17674 25050
rect 17726 24998 17738 25050
rect 17790 24998 17802 25050
rect 17854 24998 17866 25050
rect 17918 24998 22610 25050
rect 22662 24998 22674 25050
rect 22726 24998 22738 25050
rect 22790 24998 22802 25050
rect 22854 24998 22866 25050
rect 22918 24998 27610 25050
rect 27662 24998 27674 25050
rect 27726 24998 27738 25050
rect 27790 24998 27802 25050
rect 27854 24998 27866 25050
rect 27918 24998 32610 25050
rect 32662 24998 32674 25050
rect 32726 24998 32738 25050
rect 32790 24998 32802 25050
rect 32854 24998 32866 25050
rect 32918 24998 37610 25050
rect 37662 24998 37674 25050
rect 37726 24998 37738 25050
rect 37790 24998 37802 25050
rect 37854 24998 37866 25050
rect 37918 24998 38824 25050
rect 1104 24976 38824 24998
rect 1104 24506 38824 24528
rect 1104 24454 1950 24506
rect 2002 24454 2014 24506
rect 2066 24454 2078 24506
rect 2130 24454 2142 24506
rect 2194 24454 2206 24506
rect 2258 24454 6950 24506
rect 7002 24454 7014 24506
rect 7066 24454 7078 24506
rect 7130 24454 7142 24506
rect 7194 24454 7206 24506
rect 7258 24454 11950 24506
rect 12002 24454 12014 24506
rect 12066 24454 12078 24506
rect 12130 24454 12142 24506
rect 12194 24454 12206 24506
rect 12258 24454 16950 24506
rect 17002 24454 17014 24506
rect 17066 24454 17078 24506
rect 17130 24454 17142 24506
rect 17194 24454 17206 24506
rect 17258 24454 21950 24506
rect 22002 24454 22014 24506
rect 22066 24454 22078 24506
rect 22130 24454 22142 24506
rect 22194 24454 22206 24506
rect 22258 24454 26950 24506
rect 27002 24454 27014 24506
rect 27066 24454 27078 24506
rect 27130 24454 27142 24506
rect 27194 24454 27206 24506
rect 27258 24454 31950 24506
rect 32002 24454 32014 24506
rect 32066 24454 32078 24506
rect 32130 24454 32142 24506
rect 32194 24454 32206 24506
rect 32258 24454 36950 24506
rect 37002 24454 37014 24506
rect 37066 24454 37078 24506
rect 37130 24454 37142 24506
rect 37194 24454 37206 24506
rect 37258 24454 38824 24506
rect 1104 24432 38824 24454
rect 1104 23962 38824 23984
rect 1104 23910 2610 23962
rect 2662 23910 2674 23962
rect 2726 23910 2738 23962
rect 2790 23910 2802 23962
rect 2854 23910 2866 23962
rect 2918 23910 7610 23962
rect 7662 23910 7674 23962
rect 7726 23910 7738 23962
rect 7790 23910 7802 23962
rect 7854 23910 7866 23962
rect 7918 23910 12610 23962
rect 12662 23910 12674 23962
rect 12726 23910 12738 23962
rect 12790 23910 12802 23962
rect 12854 23910 12866 23962
rect 12918 23910 17610 23962
rect 17662 23910 17674 23962
rect 17726 23910 17738 23962
rect 17790 23910 17802 23962
rect 17854 23910 17866 23962
rect 17918 23910 22610 23962
rect 22662 23910 22674 23962
rect 22726 23910 22738 23962
rect 22790 23910 22802 23962
rect 22854 23910 22866 23962
rect 22918 23910 27610 23962
rect 27662 23910 27674 23962
rect 27726 23910 27738 23962
rect 27790 23910 27802 23962
rect 27854 23910 27866 23962
rect 27918 23910 32610 23962
rect 32662 23910 32674 23962
rect 32726 23910 32738 23962
rect 32790 23910 32802 23962
rect 32854 23910 32866 23962
rect 32918 23910 37610 23962
rect 37662 23910 37674 23962
rect 37726 23910 37738 23962
rect 37790 23910 37802 23962
rect 37854 23910 37866 23962
rect 37918 23910 38824 23962
rect 1104 23888 38824 23910
rect 1104 23418 38824 23440
rect 1104 23366 1950 23418
rect 2002 23366 2014 23418
rect 2066 23366 2078 23418
rect 2130 23366 2142 23418
rect 2194 23366 2206 23418
rect 2258 23366 6950 23418
rect 7002 23366 7014 23418
rect 7066 23366 7078 23418
rect 7130 23366 7142 23418
rect 7194 23366 7206 23418
rect 7258 23366 11950 23418
rect 12002 23366 12014 23418
rect 12066 23366 12078 23418
rect 12130 23366 12142 23418
rect 12194 23366 12206 23418
rect 12258 23366 16950 23418
rect 17002 23366 17014 23418
rect 17066 23366 17078 23418
rect 17130 23366 17142 23418
rect 17194 23366 17206 23418
rect 17258 23366 21950 23418
rect 22002 23366 22014 23418
rect 22066 23366 22078 23418
rect 22130 23366 22142 23418
rect 22194 23366 22206 23418
rect 22258 23366 26950 23418
rect 27002 23366 27014 23418
rect 27066 23366 27078 23418
rect 27130 23366 27142 23418
rect 27194 23366 27206 23418
rect 27258 23366 31950 23418
rect 32002 23366 32014 23418
rect 32066 23366 32078 23418
rect 32130 23366 32142 23418
rect 32194 23366 32206 23418
rect 32258 23366 36950 23418
rect 37002 23366 37014 23418
rect 37066 23366 37078 23418
rect 37130 23366 37142 23418
rect 37194 23366 37206 23418
rect 37258 23366 38824 23418
rect 1104 23344 38824 23366
rect 1104 22874 38824 22896
rect 1104 22822 2610 22874
rect 2662 22822 2674 22874
rect 2726 22822 2738 22874
rect 2790 22822 2802 22874
rect 2854 22822 2866 22874
rect 2918 22822 7610 22874
rect 7662 22822 7674 22874
rect 7726 22822 7738 22874
rect 7790 22822 7802 22874
rect 7854 22822 7866 22874
rect 7918 22822 12610 22874
rect 12662 22822 12674 22874
rect 12726 22822 12738 22874
rect 12790 22822 12802 22874
rect 12854 22822 12866 22874
rect 12918 22822 17610 22874
rect 17662 22822 17674 22874
rect 17726 22822 17738 22874
rect 17790 22822 17802 22874
rect 17854 22822 17866 22874
rect 17918 22822 22610 22874
rect 22662 22822 22674 22874
rect 22726 22822 22738 22874
rect 22790 22822 22802 22874
rect 22854 22822 22866 22874
rect 22918 22822 27610 22874
rect 27662 22822 27674 22874
rect 27726 22822 27738 22874
rect 27790 22822 27802 22874
rect 27854 22822 27866 22874
rect 27918 22822 32610 22874
rect 32662 22822 32674 22874
rect 32726 22822 32738 22874
rect 32790 22822 32802 22874
rect 32854 22822 32866 22874
rect 32918 22822 37610 22874
rect 37662 22822 37674 22874
rect 37726 22822 37738 22874
rect 37790 22822 37802 22874
rect 37854 22822 37866 22874
rect 37918 22822 38824 22874
rect 1104 22800 38824 22822
rect 1104 22330 38824 22352
rect 1104 22278 1950 22330
rect 2002 22278 2014 22330
rect 2066 22278 2078 22330
rect 2130 22278 2142 22330
rect 2194 22278 2206 22330
rect 2258 22278 6950 22330
rect 7002 22278 7014 22330
rect 7066 22278 7078 22330
rect 7130 22278 7142 22330
rect 7194 22278 7206 22330
rect 7258 22278 11950 22330
rect 12002 22278 12014 22330
rect 12066 22278 12078 22330
rect 12130 22278 12142 22330
rect 12194 22278 12206 22330
rect 12258 22278 16950 22330
rect 17002 22278 17014 22330
rect 17066 22278 17078 22330
rect 17130 22278 17142 22330
rect 17194 22278 17206 22330
rect 17258 22278 21950 22330
rect 22002 22278 22014 22330
rect 22066 22278 22078 22330
rect 22130 22278 22142 22330
rect 22194 22278 22206 22330
rect 22258 22278 26950 22330
rect 27002 22278 27014 22330
rect 27066 22278 27078 22330
rect 27130 22278 27142 22330
rect 27194 22278 27206 22330
rect 27258 22278 31950 22330
rect 32002 22278 32014 22330
rect 32066 22278 32078 22330
rect 32130 22278 32142 22330
rect 32194 22278 32206 22330
rect 32258 22278 36950 22330
rect 37002 22278 37014 22330
rect 37066 22278 37078 22330
rect 37130 22278 37142 22330
rect 37194 22278 37206 22330
rect 37258 22278 38824 22330
rect 1104 22256 38824 22278
rect 37274 21972 37280 22024
rect 37332 22012 37338 22024
rect 38289 22015 38347 22021
rect 38289 22012 38301 22015
rect 37332 21984 38301 22012
rect 37332 21972 37338 21984
rect 38289 21981 38301 21984
rect 38335 21981 38347 22015
rect 38289 21975 38347 21981
rect 38470 21836 38476 21888
rect 38528 21836 38534 21888
rect 1104 21786 38824 21808
rect 1104 21734 2610 21786
rect 2662 21734 2674 21786
rect 2726 21734 2738 21786
rect 2790 21734 2802 21786
rect 2854 21734 2866 21786
rect 2918 21734 7610 21786
rect 7662 21734 7674 21786
rect 7726 21734 7738 21786
rect 7790 21734 7802 21786
rect 7854 21734 7866 21786
rect 7918 21734 12610 21786
rect 12662 21734 12674 21786
rect 12726 21734 12738 21786
rect 12790 21734 12802 21786
rect 12854 21734 12866 21786
rect 12918 21734 17610 21786
rect 17662 21734 17674 21786
rect 17726 21734 17738 21786
rect 17790 21734 17802 21786
rect 17854 21734 17866 21786
rect 17918 21734 22610 21786
rect 22662 21734 22674 21786
rect 22726 21734 22738 21786
rect 22790 21734 22802 21786
rect 22854 21734 22866 21786
rect 22918 21734 27610 21786
rect 27662 21734 27674 21786
rect 27726 21734 27738 21786
rect 27790 21734 27802 21786
rect 27854 21734 27866 21786
rect 27918 21734 32610 21786
rect 32662 21734 32674 21786
rect 32726 21734 32738 21786
rect 32790 21734 32802 21786
rect 32854 21734 32866 21786
rect 32918 21734 37610 21786
rect 37662 21734 37674 21786
rect 37726 21734 37738 21786
rect 37790 21734 37802 21786
rect 37854 21734 37866 21786
rect 37918 21734 38824 21786
rect 1104 21712 38824 21734
rect 934 21496 940 21548
rect 992 21536 998 21548
rect 1397 21539 1455 21545
rect 1397 21536 1409 21539
rect 992 21508 1409 21536
rect 992 21496 998 21508
rect 1397 21505 1409 21508
rect 1443 21505 1455 21539
rect 1397 21499 1455 21505
rect 20438 21496 20444 21548
rect 20496 21496 20502 21548
rect 38286 21496 38292 21548
rect 38344 21496 38350 21548
rect 1578 21292 1584 21344
rect 1636 21292 1642 21344
rect 19153 21335 19211 21341
rect 19153 21301 19165 21335
rect 19199 21332 19211 21335
rect 19794 21332 19800 21344
rect 19199 21304 19800 21332
rect 19199 21301 19211 21304
rect 19153 21295 19211 21301
rect 19794 21292 19800 21304
rect 19852 21292 19858 21344
rect 38470 21292 38476 21344
rect 38528 21292 38534 21344
rect 1104 21242 38824 21264
rect 1104 21190 1950 21242
rect 2002 21190 2014 21242
rect 2066 21190 2078 21242
rect 2130 21190 2142 21242
rect 2194 21190 2206 21242
rect 2258 21190 6950 21242
rect 7002 21190 7014 21242
rect 7066 21190 7078 21242
rect 7130 21190 7142 21242
rect 7194 21190 7206 21242
rect 7258 21190 11950 21242
rect 12002 21190 12014 21242
rect 12066 21190 12078 21242
rect 12130 21190 12142 21242
rect 12194 21190 12206 21242
rect 12258 21190 16950 21242
rect 17002 21190 17014 21242
rect 17066 21190 17078 21242
rect 17130 21190 17142 21242
rect 17194 21190 17206 21242
rect 17258 21190 21950 21242
rect 22002 21190 22014 21242
rect 22066 21190 22078 21242
rect 22130 21190 22142 21242
rect 22194 21190 22206 21242
rect 22258 21190 26950 21242
rect 27002 21190 27014 21242
rect 27066 21190 27078 21242
rect 27130 21190 27142 21242
rect 27194 21190 27206 21242
rect 27258 21190 31950 21242
rect 32002 21190 32014 21242
rect 32066 21190 32078 21242
rect 32130 21190 32142 21242
rect 32194 21190 32206 21242
rect 32258 21190 36950 21242
rect 37002 21190 37014 21242
rect 37066 21190 37078 21242
rect 37130 21190 37142 21242
rect 37194 21190 37206 21242
rect 37258 21190 38824 21242
rect 1104 21168 38824 21190
rect 1578 21088 1584 21140
rect 1636 21128 1642 21140
rect 15286 21128 15292 21140
rect 1636 21100 15292 21128
rect 1636 21088 1642 21100
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 19794 20952 19800 21004
rect 19852 20952 19858 21004
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20924 1639 20927
rect 15194 20924 15200 20936
rect 1627 20896 15200 20924
rect 1627 20893 1639 20896
rect 1581 20887 1639 20893
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 19886 20884 19892 20936
rect 19944 20924 19950 20936
rect 19981 20927 20039 20933
rect 19981 20924 19993 20927
rect 19944 20896 19993 20924
rect 19944 20884 19950 20896
rect 19981 20893 19993 20896
rect 20027 20893 20039 20927
rect 19981 20887 20039 20893
rect 34514 20884 34520 20936
rect 34572 20924 34578 20936
rect 38289 20927 38347 20933
rect 38289 20924 38301 20927
rect 34572 20896 38301 20924
rect 34572 20884 34578 20896
rect 38289 20893 38301 20896
rect 38335 20893 38347 20927
rect 38289 20887 38347 20893
rect 19521 20859 19579 20865
rect 19521 20825 19533 20859
rect 19567 20856 19579 20859
rect 19702 20856 19708 20868
rect 19567 20828 19708 20856
rect 19567 20825 19579 20828
rect 19521 20819 19579 20825
rect 19702 20816 19708 20828
rect 19760 20816 19766 20868
rect 20254 20816 20260 20868
rect 20312 20816 20318 20868
rect 1394 20748 1400 20800
rect 1452 20748 1458 20800
rect 19889 20791 19947 20797
rect 19889 20757 19901 20791
rect 19935 20788 19947 20791
rect 20162 20788 20168 20800
rect 19935 20760 20168 20788
rect 19935 20757 19947 20760
rect 19889 20751 19947 20757
rect 20162 20748 20168 20760
rect 20220 20748 20226 20800
rect 38473 20791 38531 20797
rect 38473 20757 38485 20791
rect 38519 20788 38531 20791
rect 38519 20760 39068 20788
rect 38519 20757 38531 20760
rect 38473 20751 38531 20757
rect 39040 20732 39068 20760
rect 1104 20698 38824 20720
rect 1104 20646 2610 20698
rect 2662 20646 2674 20698
rect 2726 20646 2738 20698
rect 2790 20646 2802 20698
rect 2854 20646 2866 20698
rect 2918 20646 7610 20698
rect 7662 20646 7674 20698
rect 7726 20646 7738 20698
rect 7790 20646 7802 20698
rect 7854 20646 7866 20698
rect 7918 20646 12610 20698
rect 12662 20646 12674 20698
rect 12726 20646 12738 20698
rect 12790 20646 12802 20698
rect 12854 20646 12866 20698
rect 12918 20646 17610 20698
rect 17662 20646 17674 20698
rect 17726 20646 17738 20698
rect 17790 20646 17802 20698
rect 17854 20646 17866 20698
rect 17918 20646 22610 20698
rect 22662 20646 22674 20698
rect 22726 20646 22738 20698
rect 22790 20646 22802 20698
rect 22854 20646 22866 20698
rect 22918 20646 27610 20698
rect 27662 20646 27674 20698
rect 27726 20646 27738 20698
rect 27790 20646 27802 20698
rect 27854 20646 27866 20698
rect 27918 20646 32610 20698
rect 32662 20646 32674 20698
rect 32726 20646 32738 20698
rect 32790 20646 32802 20698
rect 32854 20646 32866 20698
rect 32918 20646 37610 20698
rect 37662 20646 37674 20698
rect 37726 20646 37738 20698
rect 37790 20646 37802 20698
rect 37854 20646 37866 20698
rect 37918 20646 38824 20698
rect 39022 20680 39028 20732
rect 39080 20680 39086 20732
rect 1104 20624 38824 20646
rect 15194 20544 15200 20596
rect 15252 20584 15258 20596
rect 19245 20587 19303 20593
rect 19245 20584 19257 20587
rect 15252 20556 19257 20584
rect 15252 20544 15258 20556
rect 19245 20553 19257 20556
rect 19291 20553 19303 20587
rect 19245 20547 19303 20553
rect 19794 20544 19800 20596
rect 19852 20584 19858 20596
rect 20073 20587 20131 20593
rect 20073 20584 20085 20587
rect 19852 20556 20085 20584
rect 19852 20544 19858 20556
rect 20073 20553 20085 20556
rect 20119 20553 20131 20587
rect 20073 20547 20131 20553
rect 20254 20544 20260 20596
rect 20312 20544 20318 20596
rect 20901 20587 20959 20593
rect 20901 20553 20913 20587
rect 20947 20584 20959 20587
rect 20947 20556 35894 20584
rect 20947 20553 20959 20556
rect 20901 20547 20959 20553
rect 20272 20516 20300 20544
rect 20272 20488 20484 20516
rect 19426 20408 19432 20460
rect 19484 20408 19490 20460
rect 20162 20408 20168 20460
rect 20220 20408 20226 20460
rect 20456 20457 20484 20488
rect 20257 20451 20315 20457
rect 20257 20417 20269 20451
rect 20303 20417 20315 20451
rect 20257 20411 20315 20417
rect 20441 20451 20499 20457
rect 20441 20417 20453 20451
rect 20487 20417 20499 20451
rect 20441 20411 20499 20417
rect 19518 20340 19524 20392
rect 19576 20340 19582 20392
rect 19705 20383 19763 20389
rect 19705 20349 19717 20383
rect 19751 20349 19763 20383
rect 19705 20343 19763 20349
rect 19334 20272 19340 20324
rect 19392 20312 19398 20324
rect 19720 20312 19748 20343
rect 19392 20284 19748 20312
rect 19392 20272 19398 20284
rect 19702 20204 19708 20256
rect 19760 20244 19766 20256
rect 20272 20244 20300 20411
rect 20714 20408 20720 20460
rect 20772 20408 20778 20460
rect 35866 20312 35894 20556
rect 38286 20312 38292 20324
rect 20640 20284 26234 20312
rect 35866 20284 38292 20312
rect 20640 20253 20668 20284
rect 19760 20216 20300 20244
rect 20625 20247 20683 20253
rect 19760 20204 19766 20216
rect 20625 20213 20637 20247
rect 20671 20213 20683 20247
rect 26206 20244 26234 20284
rect 38286 20272 38292 20284
rect 38344 20272 38350 20324
rect 37274 20244 37280 20256
rect 26206 20216 37280 20244
rect 20625 20207 20683 20213
rect 37274 20204 37280 20216
rect 37332 20204 37338 20256
rect 1104 20154 38824 20176
rect 1104 20102 1950 20154
rect 2002 20102 2014 20154
rect 2066 20102 2078 20154
rect 2130 20102 2142 20154
rect 2194 20102 2206 20154
rect 2258 20102 6950 20154
rect 7002 20102 7014 20154
rect 7066 20102 7078 20154
rect 7130 20102 7142 20154
rect 7194 20102 7206 20154
rect 7258 20102 11950 20154
rect 12002 20102 12014 20154
rect 12066 20102 12078 20154
rect 12130 20102 12142 20154
rect 12194 20102 12206 20154
rect 12258 20102 16950 20154
rect 17002 20102 17014 20154
rect 17066 20102 17078 20154
rect 17130 20102 17142 20154
rect 17194 20102 17206 20154
rect 17258 20102 21950 20154
rect 22002 20102 22014 20154
rect 22066 20102 22078 20154
rect 22130 20102 22142 20154
rect 22194 20102 22206 20154
rect 22258 20102 26950 20154
rect 27002 20102 27014 20154
rect 27066 20102 27078 20154
rect 27130 20102 27142 20154
rect 27194 20102 27206 20154
rect 27258 20102 31950 20154
rect 32002 20102 32014 20154
rect 32066 20102 32078 20154
rect 32130 20102 32142 20154
rect 32194 20102 32206 20154
rect 32258 20102 36950 20154
rect 37002 20102 37014 20154
rect 37066 20102 37078 20154
rect 37130 20102 37142 20154
rect 37194 20102 37206 20154
rect 37258 20102 38824 20154
rect 1104 20080 38824 20102
rect 38473 20043 38531 20049
rect 38473 20009 38485 20043
rect 38519 20040 38531 20043
rect 38519 20012 38884 20040
rect 38519 20009 38531 20012
rect 38473 20003 38531 20009
rect 38856 19984 38884 20012
rect 1581 19975 1639 19981
rect 1581 19941 1593 19975
rect 1627 19972 1639 19975
rect 19518 19972 19524 19984
rect 1627 19944 6914 19972
rect 1627 19941 1639 19944
rect 1581 19935 1639 19941
rect 6886 19904 6914 19944
rect 18340 19944 19524 19972
rect 18340 19913 18368 19944
rect 19518 19932 19524 19944
rect 19576 19972 19582 19984
rect 19886 19972 19892 19984
rect 19576 19944 19892 19972
rect 19576 19932 19582 19944
rect 19886 19932 19892 19944
rect 19944 19932 19950 19984
rect 22281 19975 22339 19981
rect 22281 19941 22293 19975
rect 22327 19972 22339 19975
rect 34514 19972 34520 19984
rect 22327 19944 34520 19972
rect 22327 19941 22339 19944
rect 22281 19935 22339 19941
rect 34514 19932 34520 19944
rect 34572 19932 34578 19984
rect 38838 19932 38844 19984
rect 38896 19932 38902 19984
rect 18325 19907 18383 19913
rect 18325 19904 18337 19907
rect 6886 19876 18337 19904
rect 18325 19873 18337 19876
rect 18371 19873 18383 19907
rect 18325 19867 18383 19873
rect 18693 19907 18751 19913
rect 18693 19873 18705 19907
rect 18739 19904 18751 19907
rect 19794 19904 19800 19916
rect 18739 19876 19800 19904
rect 18739 19873 18751 19876
rect 18693 19867 18751 19873
rect 19794 19864 19800 19876
rect 19852 19864 19858 19916
rect 934 19796 940 19848
rect 992 19836 998 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 992 19808 1409 19836
rect 992 19796 998 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 15286 19796 15292 19848
rect 15344 19836 15350 19848
rect 18785 19839 18843 19845
rect 18785 19836 18797 19839
rect 15344 19808 18797 19836
rect 15344 19796 15350 19808
rect 18785 19805 18797 19808
rect 18831 19805 18843 19839
rect 18785 19799 18843 19805
rect 19061 19839 19119 19845
rect 19061 19805 19073 19839
rect 19107 19836 19119 19839
rect 21821 19839 21879 19845
rect 21821 19836 21833 19839
rect 19107 19808 21833 19836
rect 19107 19805 19119 19808
rect 19061 19799 19119 19805
rect 21821 19805 21833 19808
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 22097 19839 22155 19845
rect 22097 19805 22109 19839
rect 22143 19836 22155 19839
rect 22278 19836 22284 19848
rect 22143 19808 22284 19836
rect 22143 19805 22155 19808
rect 22097 19799 22155 19805
rect 18800 19768 18828 19799
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 26234 19796 26240 19848
rect 26292 19836 26298 19848
rect 38289 19839 38347 19845
rect 38289 19836 38301 19839
rect 26292 19808 38301 19836
rect 26292 19796 26298 19808
rect 38289 19805 38301 19808
rect 38335 19805 38347 19839
rect 38289 19799 38347 19805
rect 19518 19768 19524 19780
rect 18800 19740 19524 19768
rect 19518 19728 19524 19740
rect 19576 19728 19582 19780
rect 21726 19728 21732 19780
rect 21784 19728 21790 19780
rect 22020 19740 26234 19768
rect 18598 19660 18604 19712
rect 18656 19700 18662 19712
rect 19702 19700 19708 19712
rect 18656 19672 19708 19700
rect 18656 19660 18662 19672
rect 19702 19660 19708 19672
rect 19760 19660 19766 19712
rect 20438 19660 20444 19712
rect 20496 19660 20502 19712
rect 22020 19709 22048 19740
rect 22005 19703 22063 19709
rect 22005 19669 22017 19703
rect 22051 19669 22063 19703
rect 26206 19700 26234 19740
rect 37274 19700 37280 19712
rect 26206 19672 37280 19700
rect 22005 19663 22063 19669
rect 37274 19660 37280 19672
rect 37332 19660 37338 19712
rect 1104 19610 38824 19632
rect 1104 19558 2610 19610
rect 2662 19558 2674 19610
rect 2726 19558 2738 19610
rect 2790 19558 2802 19610
rect 2854 19558 2866 19610
rect 2918 19558 7610 19610
rect 7662 19558 7674 19610
rect 7726 19558 7738 19610
rect 7790 19558 7802 19610
rect 7854 19558 7866 19610
rect 7918 19558 12610 19610
rect 12662 19558 12674 19610
rect 12726 19558 12738 19610
rect 12790 19558 12802 19610
rect 12854 19558 12866 19610
rect 12918 19558 17610 19610
rect 17662 19558 17674 19610
rect 17726 19558 17738 19610
rect 17790 19558 17802 19610
rect 17854 19558 17866 19610
rect 17918 19558 22610 19610
rect 22662 19558 22674 19610
rect 22726 19558 22738 19610
rect 22790 19558 22802 19610
rect 22854 19558 22866 19610
rect 22918 19558 27610 19610
rect 27662 19558 27674 19610
rect 27726 19558 27738 19610
rect 27790 19558 27802 19610
rect 27854 19558 27866 19610
rect 27918 19558 32610 19610
rect 32662 19558 32674 19610
rect 32726 19558 32738 19610
rect 32790 19558 32802 19610
rect 32854 19558 32866 19610
rect 32918 19558 37610 19610
rect 37662 19558 37674 19610
rect 37726 19558 37738 19610
rect 37790 19558 37802 19610
rect 37854 19558 37866 19610
rect 37918 19558 38824 19610
rect 1104 19536 38824 19558
rect 18966 19456 18972 19508
rect 19024 19456 19030 19508
rect 19245 19499 19303 19505
rect 19245 19465 19257 19499
rect 19291 19496 19303 19499
rect 19291 19468 21680 19496
rect 19291 19465 19303 19468
rect 19245 19459 19303 19465
rect 20993 19431 21051 19437
rect 20993 19428 21005 19431
rect 6886 19400 19656 19428
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19360 1639 19363
rect 6886 19360 6914 19400
rect 1627 19332 6914 19360
rect 18785 19363 18843 19369
rect 1627 19329 1639 19332
rect 1581 19323 1639 19329
rect 18785 19329 18797 19363
rect 18831 19360 18843 19363
rect 19061 19363 19119 19369
rect 18831 19332 19012 19360
rect 18831 19329 18843 19332
rect 18785 19323 18843 19329
rect 18984 19292 19012 19332
rect 19061 19329 19073 19363
rect 19107 19360 19119 19363
rect 19334 19360 19340 19372
rect 19107 19332 19340 19360
rect 19107 19329 19119 19332
rect 19061 19323 19119 19329
rect 19334 19320 19340 19332
rect 19392 19320 19398 19372
rect 19628 19369 19656 19400
rect 19720 19400 21005 19428
rect 19720 19372 19748 19400
rect 20993 19397 21005 19400
rect 21039 19397 21051 19431
rect 21652 19428 21680 19468
rect 21726 19456 21732 19508
rect 21784 19496 21790 19508
rect 31754 19496 31760 19508
rect 21784 19468 31760 19496
rect 21784 19456 21790 19468
rect 31754 19456 31760 19468
rect 31812 19456 31818 19508
rect 26234 19428 26240 19440
rect 21652 19400 26240 19428
rect 20993 19391 21051 19397
rect 26234 19388 26240 19400
rect 26292 19388 26298 19440
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19329 19671 19363
rect 19613 19323 19671 19329
rect 19702 19320 19708 19372
rect 19760 19320 19766 19372
rect 19886 19320 19892 19372
rect 19944 19320 19950 19372
rect 20162 19320 20168 19372
rect 20220 19320 20226 19372
rect 20625 19363 20683 19369
rect 20625 19360 20637 19363
rect 20272 19332 20637 19360
rect 20272 19292 20300 19332
rect 20625 19329 20637 19332
rect 20671 19329 20683 19363
rect 20625 19323 20683 19329
rect 21082 19320 21088 19372
rect 21140 19320 21146 19372
rect 21177 19363 21235 19369
rect 21177 19329 21189 19363
rect 21223 19329 21235 19363
rect 21177 19323 21235 19329
rect 18984 19264 20300 19292
rect 20441 19295 20499 19301
rect 20441 19261 20453 19295
rect 20487 19261 20499 19295
rect 21192 19292 21220 19323
rect 38286 19320 38292 19372
rect 38344 19320 38350 19372
rect 20441 19255 20499 19261
rect 20640 19264 21220 19292
rect 19337 19227 19395 19233
rect 19337 19193 19349 19227
rect 19383 19224 19395 19227
rect 19794 19224 19800 19236
rect 19383 19196 19800 19224
rect 19383 19193 19395 19196
rect 19337 19187 19395 19193
rect 19794 19184 19800 19196
rect 19852 19184 19858 19236
rect 1394 19116 1400 19168
rect 1452 19116 1458 19168
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 20162 19156 20168 19168
rect 19576 19128 20168 19156
rect 19576 19116 19582 19128
rect 20162 19116 20168 19128
rect 20220 19156 20226 19168
rect 20346 19156 20352 19168
rect 20220 19128 20352 19156
rect 20220 19116 20226 19128
rect 20346 19116 20352 19128
rect 20404 19156 20410 19168
rect 20456 19156 20484 19255
rect 20640 19236 20668 19264
rect 20622 19184 20628 19236
rect 20680 19184 20686 19236
rect 20404 19128 20484 19156
rect 20404 19116 20410 19128
rect 38470 19116 38476 19168
rect 38528 19116 38534 19168
rect 1104 19066 38824 19088
rect 1104 19014 1950 19066
rect 2002 19014 2014 19066
rect 2066 19014 2078 19066
rect 2130 19014 2142 19066
rect 2194 19014 2206 19066
rect 2258 19014 6950 19066
rect 7002 19014 7014 19066
rect 7066 19014 7078 19066
rect 7130 19014 7142 19066
rect 7194 19014 7206 19066
rect 7258 19014 11950 19066
rect 12002 19014 12014 19066
rect 12066 19014 12078 19066
rect 12130 19014 12142 19066
rect 12194 19014 12206 19066
rect 12258 19014 16950 19066
rect 17002 19014 17014 19066
rect 17066 19014 17078 19066
rect 17130 19014 17142 19066
rect 17194 19014 17206 19066
rect 17258 19014 21950 19066
rect 22002 19014 22014 19066
rect 22066 19014 22078 19066
rect 22130 19014 22142 19066
rect 22194 19014 22206 19066
rect 22258 19014 26950 19066
rect 27002 19014 27014 19066
rect 27066 19014 27078 19066
rect 27130 19014 27142 19066
rect 27194 19014 27206 19066
rect 27258 19014 31950 19066
rect 32002 19014 32014 19066
rect 32066 19014 32078 19066
rect 32130 19014 32142 19066
rect 32194 19014 32206 19066
rect 32258 19014 36950 19066
rect 37002 19014 37014 19066
rect 37066 19014 37078 19066
rect 37130 19014 37142 19066
rect 37194 19014 37206 19066
rect 37258 19014 38824 19066
rect 1104 18992 38824 19014
rect 20993 18955 21051 18961
rect 20993 18921 21005 18955
rect 21039 18952 21051 18955
rect 22278 18952 22284 18964
rect 21039 18924 22284 18952
rect 21039 18921 21051 18924
rect 20993 18915 21051 18921
rect 22278 18912 22284 18924
rect 22336 18912 22342 18964
rect 1581 18887 1639 18893
rect 1581 18853 1593 18887
rect 1627 18884 1639 18887
rect 18598 18884 18604 18896
rect 1627 18856 18604 18884
rect 1627 18853 1639 18856
rect 1581 18847 1639 18853
rect 18598 18844 18604 18856
rect 18656 18844 18662 18896
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 19705 18819 19763 18825
rect 19705 18816 19717 18819
rect 19484 18788 19717 18816
rect 19484 18776 19490 18788
rect 19705 18785 19717 18788
rect 19751 18785 19763 18819
rect 19705 18779 19763 18785
rect 20438 18776 20444 18828
rect 20496 18816 20502 18828
rect 20496 18788 21496 18816
rect 20496 18776 20502 18788
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 992 18720 1409 18748
rect 992 18708 998 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 19518 18708 19524 18760
rect 19576 18708 19582 18760
rect 21468 18757 21496 18788
rect 20073 18751 20131 18757
rect 20073 18717 20085 18751
rect 20119 18748 20131 18751
rect 21453 18751 21511 18757
rect 20119 18720 20852 18748
rect 20119 18717 20131 18720
rect 20073 18711 20131 18717
rect 19702 18640 19708 18692
rect 19760 18680 19766 18692
rect 20257 18683 20315 18689
rect 20257 18680 20269 18683
rect 19760 18652 20269 18680
rect 19760 18640 19766 18652
rect 20257 18649 20269 18652
rect 20303 18649 20315 18683
rect 20257 18643 20315 18649
rect 19886 18572 19892 18624
rect 19944 18612 19950 18624
rect 20165 18615 20223 18621
rect 20165 18612 20177 18615
rect 19944 18584 20177 18612
rect 19944 18572 19950 18584
rect 20165 18581 20177 18584
rect 20211 18581 20223 18615
rect 20272 18612 20300 18643
rect 20346 18640 20352 18692
rect 20404 18680 20410 18692
rect 20441 18683 20499 18689
rect 20441 18680 20453 18683
rect 20404 18652 20453 18680
rect 20404 18640 20410 18652
rect 20441 18649 20453 18652
rect 20487 18649 20499 18683
rect 20717 18683 20775 18689
rect 20717 18680 20729 18683
rect 20441 18643 20499 18649
rect 20548 18652 20729 18680
rect 20548 18612 20576 18652
rect 20717 18649 20729 18652
rect 20763 18649 20775 18683
rect 20717 18643 20775 18649
rect 20272 18584 20576 18612
rect 20165 18575 20223 18581
rect 20622 18572 20628 18624
rect 20680 18572 20686 18624
rect 20824 18621 20852 18720
rect 21453 18717 21465 18751
rect 21499 18717 21511 18751
rect 21453 18711 21511 18717
rect 37274 18708 37280 18760
rect 37332 18748 37338 18760
rect 38289 18751 38347 18757
rect 38289 18748 38301 18751
rect 37332 18720 38301 18748
rect 37332 18708 37338 18720
rect 38289 18717 38301 18720
rect 38335 18717 38347 18751
rect 38289 18711 38347 18717
rect 20809 18615 20867 18621
rect 20809 18581 20821 18615
rect 20855 18612 20867 18615
rect 21082 18612 21088 18624
rect 20855 18584 21088 18612
rect 20855 18581 20867 18584
rect 20809 18575 20867 18581
rect 21082 18572 21088 18584
rect 21140 18612 21146 18624
rect 22741 18615 22799 18621
rect 22741 18612 22753 18615
rect 21140 18584 22753 18612
rect 21140 18572 21146 18584
rect 22741 18581 22753 18584
rect 22787 18581 22799 18615
rect 22741 18575 22799 18581
rect 38470 18572 38476 18624
rect 38528 18572 38534 18624
rect 1104 18522 38824 18544
rect 1104 18470 2610 18522
rect 2662 18470 2674 18522
rect 2726 18470 2738 18522
rect 2790 18470 2802 18522
rect 2854 18470 2866 18522
rect 2918 18470 7610 18522
rect 7662 18470 7674 18522
rect 7726 18470 7738 18522
rect 7790 18470 7802 18522
rect 7854 18470 7866 18522
rect 7918 18470 12610 18522
rect 12662 18470 12674 18522
rect 12726 18470 12738 18522
rect 12790 18470 12802 18522
rect 12854 18470 12866 18522
rect 12918 18470 17610 18522
rect 17662 18470 17674 18522
rect 17726 18470 17738 18522
rect 17790 18470 17802 18522
rect 17854 18470 17866 18522
rect 17918 18470 22610 18522
rect 22662 18470 22674 18522
rect 22726 18470 22738 18522
rect 22790 18470 22802 18522
rect 22854 18470 22866 18522
rect 22918 18470 27610 18522
rect 27662 18470 27674 18522
rect 27726 18470 27738 18522
rect 27790 18470 27802 18522
rect 27854 18470 27866 18522
rect 27918 18470 32610 18522
rect 32662 18470 32674 18522
rect 32726 18470 32738 18522
rect 32790 18470 32802 18522
rect 32854 18470 32866 18522
rect 32918 18470 37610 18522
rect 37662 18470 37674 18522
rect 37726 18470 37738 18522
rect 37790 18470 37802 18522
rect 37854 18470 37866 18522
rect 37918 18470 38824 18522
rect 1104 18448 38824 18470
rect 19702 18368 19708 18420
rect 19760 18408 19766 18420
rect 19889 18411 19947 18417
rect 19889 18408 19901 18411
rect 19760 18380 19901 18408
rect 19760 18368 19766 18380
rect 19889 18377 19901 18380
rect 19935 18377 19947 18411
rect 19889 18371 19947 18377
rect 20165 18411 20223 18417
rect 20165 18377 20177 18411
rect 20211 18408 20223 18411
rect 20714 18408 20720 18420
rect 20211 18380 20720 18408
rect 20211 18377 20223 18380
rect 20165 18371 20223 18377
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 19518 18300 19524 18352
rect 19576 18300 19582 18352
rect 19981 18343 20039 18349
rect 19981 18309 19993 18343
rect 20027 18340 20039 18343
rect 21082 18340 21088 18352
rect 20027 18312 21088 18340
rect 20027 18309 20039 18312
rect 19981 18303 20039 18309
rect 21082 18300 21088 18312
rect 21140 18300 21146 18352
rect 19797 18275 19855 18281
rect 19797 18241 19809 18275
rect 19843 18272 19855 18275
rect 19886 18272 19892 18284
rect 19843 18244 19892 18272
rect 19843 18241 19855 18244
rect 19797 18235 19855 18241
rect 19886 18232 19892 18244
rect 19944 18272 19950 18284
rect 20622 18272 20628 18284
rect 19944 18244 20628 18272
rect 19944 18232 19950 18244
rect 20622 18232 20628 18244
rect 20680 18232 20686 18284
rect 1104 17978 38824 18000
rect 1104 17926 1950 17978
rect 2002 17926 2014 17978
rect 2066 17926 2078 17978
rect 2130 17926 2142 17978
rect 2194 17926 2206 17978
rect 2258 17926 6950 17978
rect 7002 17926 7014 17978
rect 7066 17926 7078 17978
rect 7130 17926 7142 17978
rect 7194 17926 7206 17978
rect 7258 17926 11950 17978
rect 12002 17926 12014 17978
rect 12066 17926 12078 17978
rect 12130 17926 12142 17978
rect 12194 17926 12206 17978
rect 12258 17926 16950 17978
rect 17002 17926 17014 17978
rect 17066 17926 17078 17978
rect 17130 17926 17142 17978
rect 17194 17926 17206 17978
rect 17258 17926 21950 17978
rect 22002 17926 22014 17978
rect 22066 17926 22078 17978
rect 22130 17926 22142 17978
rect 22194 17926 22206 17978
rect 22258 17926 26950 17978
rect 27002 17926 27014 17978
rect 27066 17926 27078 17978
rect 27130 17926 27142 17978
rect 27194 17926 27206 17978
rect 27258 17926 31950 17978
rect 32002 17926 32014 17978
rect 32066 17926 32078 17978
rect 32130 17926 32142 17978
rect 32194 17926 32206 17978
rect 32258 17926 36950 17978
rect 37002 17926 37014 17978
rect 37066 17926 37078 17978
rect 37130 17926 37142 17978
rect 37194 17926 37206 17978
rect 37258 17926 38824 17978
rect 1104 17904 38824 17926
rect 31754 17824 31760 17876
rect 31812 17864 31818 17876
rect 34514 17864 34520 17876
rect 31812 17836 34520 17864
rect 31812 17824 31818 17836
rect 34514 17824 34520 17836
rect 34572 17824 34578 17876
rect 1104 17434 38824 17456
rect 1104 17382 2610 17434
rect 2662 17382 2674 17434
rect 2726 17382 2738 17434
rect 2790 17382 2802 17434
rect 2854 17382 2866 17434
rect 2918 17382 7610 17434
rect 7662 17382 7674 17434
rect 7726 17382 7738 17434
rect 7790 17382 7802 17434
rect 7854 17382 7866 17434
rect 7918 17382 12610 17434
rect 12662 17382 12674 17434
rect 12726 17382 12738 17434
rect 12790 17382 12802 17434
rect 12854 17382 12866 17434
rect 12918 17382 17610 17434
rect 17662 17382 17674 17434
rect 17726 17382 17738 17434
rect 17790 17382 17802 17434
rect 17854 17382 17866 17434
rect 17918 17382 22610 17434
rect 22662 17382 22674 17434
rect 22726 17382 22738 17434
rect 22790 17382 22802 17434
rect 22854 17382 22866 17434
rect 22918 17382 27610 17434
rect 27662 17382 27674 17434
rect 27726 17382 27738 17434
rect 27790 17382 27802 17434
rect 27854 17382 27866 17434
rect 27918 17382 32610 17434
rect 32662 17382 32674 17434
rect 32726 17382 32738 17434
rect 32790 17382 32802 17434
rect 32854 17382 32866 17434
rect 32918 17382 37610 17434
rect 37662 17382 37674 17434
rect 37726 17382 37738 17434
rect 37790 17382 37802 17434
rect 37854 17382 37866 17434
rect 37918 17382 38824 17434
rect 1104 17360 38824 17382
rect 1104 16890 38824 16912
rect 1104 16838 1950 16890
rect 2002 16838 2014 16890
rect 2066 16838 2078 16890
rect 2130 16838 2142 16890
rect 2194 16838 2206 16890
rect 2258 16838 6950 16890
rect 7002 16838 7014 16890
rect 7066 16838 7078 16890
rect 7130 16838 7142 16890
rect 7194 16838 7206 16890
rect 7258 16838 11950 16890
rect 12002 16838 12014 16890
rect 12066 16838 12078 16890
rect 12130 16838 12142 16890
rect 12194 16838 12206 16890
rect 12258 16838 16950 16890
rect 17002 16838 17014 16890
rect 17066 16838 17078 16890
rect 17130 16838 17142 16890
rect 17194 16838 17206 16890
rect 17258 16838 21950 16890
rect 22002 16838 22014 16890
rect 22066 16838 22078 16890
rect 22130 16838 22142 16890
rect 22194 16838 22206 16890
rect 22258 16838 26950 16890
rect 27002 16838 27014 16890
rect 27066 16838 27078 16890
rect 27130 16838 27142 16890
rect 27194 16838 27206 16890
rect 27258 16838 31950 16890
rect 32002 16838 32014 16890
rect 32066 16838 32078 16890
rect 32130 16838 32142 16890
rect 32194 16838 32206 16890
rect 32258 16838 36950 16890
rect 37002 16838 37014 16890
rect 37066 16838 37078 16890
rect 37130 16838 37142 16890
rect 37194 16838 37206 16890
rect 37258 16838 38824 16890
rect 1104 16816 38824 16838
rect 1104 16346 38824 16368
rect 1104 16294 2610 16346
rect 2662 16294 2674 16346
rect 2726 16294 2738 16346
rect 2790 16294 2802 16346
rect 2854 16294 2866 16346
rect 2918 16294 7610 16346
rect 7662 16294 7674 16346
rect 7726 16294 7738 16346
rect 7790 16294 7802 16346
rect 7854 16294 7866 16346
rect 7918 16294 12610 16346
rect 12662 16294 12674 16346
rect 12726 16294 12738 16346
rect 12790 16294 12802 16346
rect 12854 16294 12866 16346
rect 12918 16294 17610 16346
rect 17662 16294 17674 16346
rect 17726 16294 17738 16346
rect 17790 16294 17802 16346
rect 17854 16294 17866 16346
rect 17918 16294 22610 16346
rect 22662 16294 22674 16346
rect 22726 16294 22738 16346
rect 22790 16294 22802 16346
rect 22854 16294 22866 16346
rect 22918 16294 27610 16346
rect 27662 16294 27674 16346
rect 27726 16294 27738 16346
rect 27790 16294 27802 16346
rect 27854 16294 27866 16346
rect 27918 16294 32610 16346
rect 32662 16294 32674 16346
rect 32726 16294 32738 16346
rect 32790 16294 32802 16346
rect 32854 16294 32866 16346
rect 32918 16294 37610 16346
rect 37662 16294 37674 16346
rect 37726 16294 37738 16346
rect 37790 16294 37802 16346
rect 37854 16294 37866 16346
rect 37918 16294 38824 16346
rect 1104 16272 38824 16294
rect 1104 15802 38824 15824
rect 1104 15750 1950 15802
rect 2002 15750 2014 15802
rect 2066 15750 2078 15802
rect 2130 15750 2142 15802
rect 2194 15750 2206 15802
rect 2258 15750 6950 15802
rect 7002 15750 7014 15802
rect 7066 15750 7078 15802
rect 7130 15750 7142 15802
rect 7194 15750 7206 15802
rect 7258 15750 11950 15802
rect 12002 15750 12014 15802
rect 12066 15750 12078 15802
rect 12130 15750 12142 15802
rect 12194 15750 12206 15802
rect 12258 15750 16950 15802
rect 17002 15750 17014 15802
rect 17066 15750 17078 15802
rect 17130 15750 17142 15802
rect 17194 15750 17206 15802
rect 17258 15750 21950 15802
rect 22002 15750 22014 15802
rect 22066 15750 22078 15802
rect 22130 15750 22142 15802
rect 22194 15750 22206 15802
rect 22258 15750 26950 15802
rect 27002 15750 27014 15802
rect 27066 15750 27078 15802
rect 27130 15750 27142 15802
rect 27194 15750 27206 15802
rect 27258 15750 31950 15802
rect 32002 15750 32014 15802
rect 32066 15750 32078 15802
rect 32130 15750 32142 15802
rect 32194 15750 32206 15802
rect 32258 15750 36950 15802
rect 37002 15750 37014 15802
rect 37066 15750 37078 15802
rect 37130 15750 37142 15802
rect 37194 15750 37206 15802
rect 37258 15750 38824 15802
rect 1104 15728 38824 15750
rect 1104 15258 38824 15280
rect 1104 15206 2610 15258
rect 2662 15206 2674 15258
rect 2726 15206 2738 15258
rect 2790 15206 2802 15258
rect 2854 15206 2866 15258
rect 2918 15206 7610 15258
rect 7662 15206 7674 15258
rect 7726 15206 7738 15258
rect 7790 15206 7802 15258
rect 7854 15206 7866 15258
rect 7918 15206 12610 15258
rect 12662 15206 12674 15258
rect 12726 15206 12738 15258
rect 12790 15206 12802 15258
rect 12854 15206 12866 15258
rect 12918 15206 17610 15258
rect 17662 15206 17674 15258
rect 17726 15206 17738 15258
rect 17790 15206 17802 15258
rect 17854 15206 17866 15258
rect 17918 15206 22610 15258
rect 22662 15206 22674 15258
rect 22726 15206 22738 15258
rect 22790 15206 22802 15258
rect 22854 15206 22866 15258
rect 22918 15206 27610 15258
rect 27662 15206 27674 15258
rect 27726 15206 27738 15258
rect 27790 15206 27802 15258
rect 27854 15206 27866 15258
rect 27918 15206 32610 15258
rect 32662 15206 32674 15258
rect 32726 15206 32738 15258
rect 32790 15206 32802 15258
rect 32854 15206 32866 15258
rect 32918 15206 37610 15258
rect 37662 15206 37674 15258
rect 37726 15206 37738 15258
rect 37790 15206 37802 15258
rect 37854 15206 37866 15258
rect 37918 15206 38824 15258
rect 1104 15184 38824 15206
rect 1104 14714 38824 14736
rect 1104 14662 1950 14714
rect 2002 14662 2014 14714
rect 2066 14662 2078 14714
rect 2130 14662 2142 14714
rect 2194 14662 2206 14714
rect 2258 14662 6950 14714
rect 7002 14662 7014 14714
rect 7066 14662 7078 14714
rect 7130 14662 7142 14714
rect 7194 14662 7206 14714
rect 7258 14662 11950 14714
rect 12002 14662 12014 14714
rect 12066 14662 12078 14714
rect 12130 14662 12142 14714
rect 12194 14662 12206 14714
rect 12258 14662 16950 14714
rect 17002 14662 17014 14714
rect 17066 14662 17078 14714
rect 17130 14662 17142 14714
rect 17194 14662 17206 14714
rect 17258 14662 21950 14714
rect 22002 14662 22014 14714
rect 22066 14662 22078 14714
rect 22130 14662 22142 14714
rect 22194 14662 22206 14714
rect 22258 14662 26950 14714
rect 27002 14662 27014 14714
rect 27066 14662 27078 14714
rect 27130 14662 27142 14714
rect 27194 14662 27206 14714
rect 27258 14662 31950 14714
rect 32002 14662 32014 14714
rect 32066 14662 32078 14714
rect 32130 14662 32142 14714
rect 32194 14662 32206 14714
rect 32258 14662 36950 14714
rect 37002 14662 37014 14714
rect 37066 14662 37078 14714
rect 37130 14662 37142 14714
rect 37194 14662 37206 14714
rect 37258 14662 38824 14714
rect 1104 14640 38824 14662
rect 1104 14170 38824 14192
rect 1104 14118 2610 14170
rect 2662 14118 2674 14170
rect 2726 14118 2738 14170
rect 2790 14118 2802 14170
rect 2854 14118 2866 14170
rect 2918 14118 7610 14170
rect 7662 14118 7674 14170
rect 7726 14118 7738 14170
rect 7790 14118 7802 14170
rect 7854 14118 7866 14170
rect 7918 14118 12610 14170
rect 12662 14118 12674 14170
rect 12726 14118 12738 14170
rect 12790 14118 12802 14170
rect 12854 14118 12866 14170
rect 12918 14118 17610 14170
rect 17662 14118 17674 14170
rect 17726 14118 17738 14170
rect 17790 14118 17802 14170
rect 17854 14118 17866 14170
rect 17918 14118 22610 14170
rect 22662 14118 22674 14170
rect 22726 14118 22738 14170
rect 22790 14118 22802 14170
rect 22854 14118 22866 14170
rect 22918 14118 27610 14170
rect 27662 14118 27674 14170
rect 27726 14118 27738 14170
rect 27790 14118 27802 14170
rect 27854 14118 27866 14170
rect 27918 14118 32610 14170
rect 32662 14118 32674 14170
rect 32726 14118 32738 14170
rect 32790 14118 32802 14170
rect 32854 14118 32866 14170
rect 32918 14118 37610 14170
rect 37662 14118 37674 14170
rect 37726 14118 37738 14170
rect 37790 14118 37802 14170
rect 37854 14118 37866 14170
rect 37918 14118 38824 14170
rect 1104 14096 38824 14118
rect 1104 13626 38824 13648
rect 1104 13574 1950 13626
rect 2002 13574 2014 13626
rect 2066 13574 2078 13626
rect 2130 13574 2142 13626
rect 2194 13574 2206 13626
rect 2258 13574 6950 13626
rect 7002 13574 7014 13626
rect 7066 13574 7078 13626
rect 7130 13574 7142 13626
rect 7194 13574 7206 13626
rect 7258 13574 11950 13626
rect 12002 13574 12014 13626
rect 12066 13574 12078 13626
rect 12130 13574 12142 13626
rect 12194 13574 12206 13626
rect 12258 13574 16950 13626
rect 17002 13574 17014 13626
rect 17066 13574 17078 13626
rect 17130 13574 17142 13626
rect 17194 13574 17206 13626
rect 17258 13574 21950 13626
rect 22002 13574 22014 13626
rect 22066 13574 22078 13626
rect 22130 13574 22142 13626
rect 22194 13574 22206 13626
rect 22258 13574 26950 13626
rect 27002 13574 27014 13626
rect 27066 13574 27078 13626
rect 27130 13574 27142 13626
rect 27194 13574 27206 13626
rect 27258 13574 31950 13626
rect 32002 13574 32014 13626
rect 32066 13574 32078 13626
rect 32130 13574 32142 13626
rect 32194 13574 32206 13626
rect 32258 13574 36950 13626
rect 37002 13574 37014 13626
rect 37066 13574 37078 13626
rect 37130 13574 37142 13626
rect 37194 13574 37206 13626
rect 37258 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 2610 13082
rect 2662 13030 2674 13082
rect 2726 13030 2738 13082
rect 2790 13030 2802 13082
rect 2854 13030 2866 13082
rect 2918 13030 7610 13082
rect 7662 13030 7674 13082
rect 7726 13030 7738 13082
rect 7790 13030 7802 13082
rect 7854 13030 7866 13082
rect 7918 13030 12610 13082
rect 12662 13030 12674 13082
rect 12726 13030 12738 13082
rect 12790 13030 12802 13082
rect 12854 13030 12866 13082
rect 12918 13030 17610 13082
rect 17662 13030 17674 13082
rect 17726 13030 17738 13082
rect 17790 13030 17802 13082
rect 17854 13030 17866 13082
rect 17918 13030 22610 13082
rect 22662 13030 22674 13082
rect 22726 13030 22738 13082
rect 22790 13030 22802 13082
rect 22854 13030 22866 13082
rect 22918 13030 27610 13082
rect 27662 13030 27674 13082
rect 27726 13030 27738 13082
rect 27790 13030 27802 13082
rect 27854 13030 27866 13082
rect 27918 13030 32610 13082
rect 32662 13030 32674 13082
rect 32726 13030 32738 13082
rect 32790 13030 32802 13082
rect 32854 13030 32866 13082
rect 32918 13030 37610 13082
rect 37662 13030 37674 13082
rect 37726 13030 37738 13082
rect 37790 13030 37802 13082
rect 37854 13030 37866 13082
rect 37918 13030 38824 13082
rect 1104 13008 38824 13030
rect 1104 12538 38824 12560
rect 1104 12486 1950 12538
rect 2002 12486 2014 12538
rect 2066 12486 2078 12538
rect 2130 12486 2142 12538
rect 2194 12486 2206 12538
rect 2258 12486 6950 12538
rect 7002 12486 7014 12538
rect 7066 12486 7078 12538
rect 7130 12486 7142 12538
rect 7194 12486 7206 12538
rect 7258 12486 11950 12538
rect 12002 12486 12014 12538
rect 12066 12486 12078 12538
rect 12130 12486 12142 12538
rect 12194 12486 12206 12538
rect 12258 12486 16950 12538
rect 17002 12486 17014 12538
rect 17066 12486 17078 12538
rect 17130 12486 17142 12538
rect 17194 12486 17206 12538
rect 17258 12486 21950 12538
rect 22002 12486 22014 12538
rect 22066 12486 22078 12538
rect 22130 12486 22142 12538
rect 22194 12486 22206 12538
rect 22258 12486 26950 12538
rect 27002 12486 27014 12538
rect 27066 12486 27078 12538
rect 27130 12486 27142 12538
rect 27194 12486 27206 12538
rect 27258 12486 31950 12538
rect 32002 12486 32014 12538
rect 32066 12486 32078 12538
rect 32130 12486 32142 12538
rect 32194 12486 32206 12538
rect 32258 12486 36950 12538
rect 37002 12486 37014 12538
rect 37066 12486 37078 12538
rect 37130 12486 37142 12538
rect 37194 12486 37206 12538
rect 37258 12486 38824 12538
rect 1104 12464 38824 12486
rect 1104 11994 38824 12016
rect 1104 11942 2610 11994
rect 2662 11942 2674 11994
rect 2726 11942 2738 11994
rect 2790 11942 2802 11994
rect 2854 11942 2866 11994
rect 2918 11942 7610 11994
rect 7662 11942 7674 11994
rect 7726 11942 7738 11994
rect 7790 11942 7802 11994
rect 7854 11942 7866 11994
rect 7918 11942 12610 11994
rect 12662 11942 12674 11994
rect 12726 11942 12738 11994
rect 12790 11942 12802 11994
rect 12854 11942 12866 11994
rect 12918 11942 17610 11994
rect 17662 11942 17674 11994
rect 17726 11942 17738 11994
rect 17790 11942 17802 11994
rect 17854 11942 17866 11994
rect 17918 11942 22610 11994
rect 22662 11942 22674 11994
rect 22726 11942 22738 11994
rect 22790 11942 22802 11994
rect 22854 11942 22866 11994
rect 22918 11942 27610 11994
rect 27662 11942 27674 11994
rect 27726 11942 27738 11994
rect 27790 11942 27802 11994
rect 27854 11942 27866 11994
rect 27918 11942 32610 11994
rect 32662 11942 32674 11994
rect 32726 11942 32738 11994
rect 32790 11942 32802 11994
rect 32854 11942 32866 11994
rect 32918 11942 37610 11994
rect 37662 11942 37674 11994
rect 37726 11942 37738 11994
rect 37790 11942 37802 11994
rect 37854 11942 37866 11994
rect 37918 11942 38824 11994
rect 1104 11920 38824 11942
rect 1104 11450 38824 11472
rect 1104 11398 1950 11450
rect 2002 11398 2014 11450
rect 2066 11398 2078 11450
rect 2130 11398 2142 11450
rect 2194 11398 2206 11450
rect 2258 11398 6950 11450
rect 7002 11398 7014 11450
rect 7066 11398 7078 11450
rect 7130 11398 7142 11450
rect 7194 11398 7206 11450
rect 7258 11398 11950 11450
rect 12002 11398 12014 11450
rect 12066 11398 12078 11450
rect 12130 11398 12142 11450
rect 12194 11398 12206 11450
rect 12258 11398 16950 11450
rect 17002 11398 17014 11450
rect 17066 11398 17078 11450
rect 17130 11398 17142 11450
rect 17194 11398 17206 11450
rect 17258 11398 21950 11450
rect 22002 11398 22014 11450
rect 22066 11398 22078 11450
rect 22130 11398 22142 11450
rect 22194 11398 22206 11450
rect 22258 11398 26950 11450
rect 27002 11398 27014 11450
rect 27066 11398 27078 11450
rect 27130 11398 27142 11450
rect 27194 11398 27206 11450
rect 27258 11398 31950 11450
rect 32002 11398 32014 11450
rect 32066 11398 32078 11450
rect 32130 11398 32142 11450
rect 32194 11398 32206 11450
rect 32258 11398 36950 11450
rect 37002 11398 37014 11450
rect 37066 11398 37078 11450
rect 37130 11398 37142 11450
rect 37194 11398 37206 11450
rect 37258 11398 38824 11450
rect 1104 11376 38824 11398
rect 1104 10906 38824 10928
rect 1104 10854 2610 10906
rect 2662 10854 2674 10906
rect 2726 10854 2738 10906
rect 2790 10854 2802 10906
rect 2854 10854 2866 10906
rect 2918 10854 7610 10906
rect 7662 10854 7674 10906
rect 7726 10854 7738 10906
rect 7790 10854 7802 10906
rect 7854 10854 7866 10906
rect 7918 10854 12610 10906
rect 12662 10854 12674 10906
rect 12726 10854 12738 10906
rect 12790 10854 12802 10906
rect 12854 10854 12866 10906
rect 12918 10854 17610 10906
rect 17662 10854 17674 10906
rect 17726 10854 17738 10906
rect 17790 10854 17802 10906
rect 17854 10854 17866 10906
rect 17918 10854 22610 10906
rect 22662 10854 22674 10906
rect 22726 10854 22738 10906
rect 22790 10854 22802 10906
rect 22854 10854 22866 10906
rect 22918 10854 27610 10906
rect 27662 10854 27674 10906
rect 27726 10854 27738 10906
rect 27790 10854 27802 10906
rect 27854 10854 27866 10906
rect 27918 10854 32610 10906
rect 32662 10854 32674 10906
rect 32726 10854 32738 10906
rect 32790 10854 32802 10906
rect 32854 10854 32866 10906
rect 32918 10854 37610 10906
rect 37662 10854 37674 10906
rect 37726 10854 37738 10906
rect 37790 10854 37802 10906
rect 37854 10854 37866 10906
rect 37918 10854 38824 10906
rect 1104 10832 38824 10854
rect 1104 10362 38824 10384
rect 1104 10310 1950 10362
rect 2002 10310 2014 10362
rect 2066 10310 2078 10362
rect 2130 10310 2142 10362
rect 2194 10310 2206 10362
rect 2258 10310 6950 10362
rect 7002 10310 7014 10362
rect 7066 10310 7078 10362
rect 7130 10310 7142 10362
rect 7194 10310 7206 10362
rect 7258 10310 11950 10362
rect 12002 10310 12014 10362
rect 12066 10310 12078 10362
rect 12130 10310 12142 10362
rect 12194 10310 12206 10362
rect 12258 10310 16950 10362
rect 17002 10310 17014 10362
rect 17066 10310 17078 10362
rect 17130 10310 17142 10362
rect 17194 10310 17206 10362
rect 17258 10310 21950 10362
rect 22002 10310 22014 10362
rect 22066 10310 22078 10362
rect 22130 10310 22142 10362
rect 22194 10310 22206 10362
rect 22258 10310 26950 10362
rect 27002 10310 27014 10362
rect 27066 10310 27078 10362
rect 27130 10310 27142 10362
rect 27194 10310 27206 10362
rect 27258 10310 31950 10362
rect 32002 10310 32014 10362
rect 32066 10310 32078 10362
rect 32130 10310 32142 10362
rect 32194 10310 32206 10362
rect 32258 10310 36950 10362
rect 37002 10310 37014 10362
rect 37066 10310 37078 10362
rect 37130 10310 37142 10362
rect 37194 10310 37206 10362
rect 37258 10310 38824 10362
rect 1104 10288 38824 10310
rect 1104 9818 38824 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 7610 9818
rect 7662 9766 7674 9818
rect 7726 9766 7738 9818
rect 7790 9766 7802 9818
rect 7854 9766 7866 9818
rect 7918 9766 12610 9818
rect 12662 9766 12674 9818
rect 12726 9766 12738 9818
rect 12790 9766 12802 9818
rect 12854 9766 12866 9818
rect 12918 9766 17610 9818
rect 17662 9766 17674 9818
rect 17726 9766 17738 9818
rect 17790 9766 17802 9818
rect 17854 9766 17866 9818
rect 17918 9766 22610 9818
rect 22662 9766 22674 9818
rect 22726 9766 22738 9818
rect 22790 9766 22802 9818
rect 22854 9766 22866 9818
rect 22918 9766 27610 9818
rect 27662 9766 27674 9818
rect 27726 9766 27738 9818
rect 27790 9766 27802 9818
rect 27854 9766 27866 9818
rect 27918 9766 32610 9818
rect 32662 9766 32674 9818
rect 32726 9766 32738 9818
rect 32790 9766 32802 9818
rect 32854 9766 32866 9818
rect 32918 9766 37610 9818
rect 37662 9766 37674 9818
rect 37726 9766 37738 9818
rect 37790 9766 37802 9818
rect 37854 9766 37866 9818
rect 37918 9766 38824 9818
rect 1104 9744 38824 9766
rect 1104 9274 38824 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 6950 9274
rect 7002 9222 7014 9274
rect 7066 9222 7078 9274
rect 7130 9222 7142 9274
rect 7194 9222 7206 9274
rect 7258 9222 11950 9274
rect 12002 9222 12014 9274
rect 12066 9222 12078 9274
rect 12130 9222 12142 9274
rect 12194 9222 12206 9274
rect 12258 9222 16950 9274
rect 17002 9222 17014 9274
rect 17066 9222 17078 9274
rect 17130 9222 17142 9274
rect 17194 9222 17206 9274
rect 17258 9222 21950 9274
rect 22002 9222 22014 9274
rect 22066 9222 22078 9274
rect 22130 9222 22142 9274
rect 22194 9222 22206 9274
rect 22258 9222 26950 9274
rect 27002 9222 27014 9274
rect 27066 9222 27078 9274
rect 27130 9222 27142 9274
rect 27194 9222 27206 9274
rect 27258 9222 31950 9274
rect 32002 9222 32014 9274
rect 32066 9222 32078 9274
rect 32130 9222 32142 9274
rect 32194 9222 32206 9274
rect 32258 9222 36950 9274
rect 37002 9222 37014 9274
rect 37066 9222 37078 9274
rect 37130 9222 37142 9274
rect 37194 9222 37206 9274
rect 37258 9222 38824 9274
rect 1104 9200 38824 9222
rect 1104 8730 38824 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 7610 8730
rect 7662 8678 7674 8730
rect 7726 8678 7738 8730
rect 7790 8678 7802 8730
rect 7854 8678 7866 8730
rect 7918 8678 12610 8730
rect 12662 8678 12674 8730
rect 12726 8678 12738 8730
rect 12790 8678 12802 8730
rect 12854 8678 12866 8730
rect 12918 8678 17610 8730
rect 17662 8678 17674 8730
rect 17726 8678 17738 8730
rect 17790 8678 17802 8730
rect 17854 8678 17866 8730
rect 17918 8678 22610 8730
rect 22662 8678 22674 8730
rect 22726 8678 22738 8730
rect 22790 8678 22802 8730
rect 22854 8678 22866 8730
rect 22918 8678 27610 8730
rect 27662 8678 27674 8730
rect 27726 8678 27738 8730
rect 27790 8678 27802 8730
rect 27854 8678 27866 8730
rect 27918 8678 32610 8730
rect 32662 8678 32674 8730
rect 32726 8678 32738 8730
rect 32790 8678 32802 8730
rect 32854 8678 32866 8730
rect 32918 8678 37610 8730
rect 37662 8678 37674 8730
rect 37726 8678 37738 8730
rect 37790 8678 37802 8730
rect 37854 8678 37866 8730
rect 37918 8678 38824 8730
rect 1104 8656 38824 8678
rect 1104 8186 38824 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 6950 8186
rect 7002 8134 7014 8186
rect 7066 8134 7078 8186
rect 7130 8134 7142 8186
rect 7194 8134 7206 8186
rect 7258 8134 11950 8186
rect 12002 8134 12014 8186
rect 12066 8134 12078 8186
rect 12130 8134 12142 8186
rect 12194 8134 12206 8186
rect 12258 8134 16950 8186
rect 17002 8134 17014 8186
rect 17066 8134 17078 8186
rect 17130 8134 17142 8186
rect 17194 8134 17206 8186
rect 17258 8134 21950 8186
rect 22002 8134 22014 8186
rect 22066 8134 22078 8186
rect 22130 8134 22142 8186
rect 22194 8134 22206 8186
rect 22258 8134 26950 8186
rect 27002 8134 27014 8186
rect 27066 8134 27078 8186
rect 27130 8134 27142 8186
rect 27194 8134 27206 8186
rect 27258 8134 31950 8186
rect 32002 8134 32014 8186
rect 32066 8134 32078 8186
rect 32130 8134 32142 8186
rect 32194 8134 32206 8186
rect 32258 8134 36950 8186
rect 37002 8134 37014 8186
rect 37066 8134 37078 8186
rect 37130 8134 37142 8186
rect 37194 8134 37206 8186
rect 37258 8134 38824 8186
rect 1104 8112 38824 8134
rect 1104 7642 38824 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 7610 7642
rect 7662 7590 7674 7642
rect 7726 7590 7738 7642
rect 7790 7590 7802 7642
rect 7854 7590 7866 7642
rect 7918 7590 12610 7642
rect 12662 7590 12674 7642
rect 12726 7590 12738 7642
rect 12790 7590 12802 7642
rect 12854 7590 12866 7642
rect 12918 7590 17610 7642
rect 17662 7590 17674 7642
rect 17726 7590 17738 7642
rect 17790 7590 17802 7642
rect 17854 7590 17866 7642
rect 17918 7590 22610 7642
rect 22662 7590 22674 7642
rect 22726 7590 22738 7642
rect 22790 7590 22802 7642
rect 22854 7590 22866 7642
rect 22918 7590 27610 7642
rect 27662 7590 27674 7642
rect 27726 7590 27738 7642
rect 27790 7590 27802 7642
rect 27854 7590 27866 7642
rect 27918 7590 32610 7642
rect 32662 7590 32674 7642
rect 32726 7590 32738 7642
rect 32790 7590 32802 7642
rect 32854 7590 32866 7642
rect 32918 7590 37610 7642
rect 37662 7590 37674 7642
rect 37726 7590 37738 7642
rect 37790 7590 37802 7642
rect 37854 7590 37866 7642
rect 37918 7590 38824 7642
rect 1104 7568 38824 7590
rect 1104 7098 38824 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 6950 7098
rect 7002 7046 7014 7098
rect 7066 7046 7078 7098
rect 7130 7046 7142 7098
rect 7194 7046 7206 7098
rect 7258 7046 11950 7098
rect 12002 7046 12014 7098
rect 12066 7046 12078 7098
rect 12130 7046 12142 7098
rect 12194 7046 12206 7098
rect 12258 7046 16950 7098
rect 17002 7046 17014 7098
rect 17066 7046 17078 7098
rect 17130 7046 17142 7098
rect 17194 7046 17206 7098
rect 17258 7046 21950 7098
rect 22002 7046 22014 7098
rect 22066 7046 22078 7098
rect 22130 7046 22142 7098
rect 22194 7046 22206 7098
rect 22258 7046 26950 7098
rect 27002 7046 27014 7098
rect 27066 7046 27078 7098
rect 27130 7046 27142 7098
rect 27194 7046 27206 7098
rect 27258 7046 31950 7098
rect 32002 7046 32014 7098
rect 32066 7046 32078 7098
rect 32130 7046 32142 7098
rect 32194 7046 32206 7098
rect 32258 7046 36950 7098
rect 37002 7046 37014 7098
rect 37066 7046 37078 7098
rect 37130 7046 37142 7098
rect 37194 7046 37206 7098
rect 37258 7046 38824 7098
rect 1104 7024 38824 7046
rect 1104 6554 38824 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 7610 6554
rect 7662 6502 7674 6554
rect 7726 6502 7738 6554
rect 7790 6502 7802 6554
rect 7854 6502 7866 6554
rect 7918 6502 12610 6554
rect 12662 6502 12674 6554
rect 12726 6502 12738 6554
rect 12790 6502 12802 6554
rect 12854 6502 12866 6554
rect 12918 6502 17610 6554
rect 17662 6502 17674 6554
rect 17726 6502 17738 6554
rect 17790 6502 17802 6554
rect 17854 6502 17866 6554
rect 17918 6502 22610 6554
rect 22662 6502 22674 6554
rect 22726 6502 22738 6554
rect 22790 6502 22802 6554
rect 22854 6502 22866 6554
rect 22918 6502 27610 6554
rect 27662 6502 27674 6554
rect 27726 6502 27738 6554
rect 27790 6502 27802 6554
rect 27854 6502 27866 6554
rect 27918 6502 32610 6554
rect 32662 6502 32674 6554
rect 32726 6502 32738 6554
rect 32790 6502 32802 6554
rect 32854 6502 32866 6554
rect 32918 6502 37610 6554
rect 37662 6502 37674 6554
rect 37726 6502 37738 6554
rect 37790 6502 37802 6554
rect 37854 6502 37866 6554
rect 37918 6502 38824 6554
rect 1104 6480 38824 6502
rect 1104 6010 38824 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 6950 6010
rect 7002 5958 7014 6010
rect 7066 5958 7078 6010
rect 7130 5958 7142 6010
rect 7194 5958 7206 6010
rect 7258 5958 11950 6010
rect 12002 5958 12014 6010
rect 12066 5958 12078 6010
rect 12130 5958 12142 6010
rect 12194 5958 12206 6010
rect 12258 5958 16950 6010
rect 17002 5958 17014 6010
rect 17066 5958 17078 6010
rect 17130 5958 17142 6010
rect 17194 5958 17206 6010
rect 17258 5958 21950 6010
rect 22002 5958 22014 6010
rect 22066 5958 22078 6010
rect 22130 5958 22142 6010
rect 22194 5958 22206 6010
rect 22258 5958 26950 6010
rect 27002 5958 27014 6010
rect 27066 5958 27078 6010
rect 27130 5958 27142 6010
rect 27194 5958 27206 6010
rect 27258 5958 31950 6010
rect 32002 5958 32014 6010
rect 32066 5958 32078 6010
rect 32130 5958 32142 6010
rect 32194 5958 32206 6010
rect 32258 5958 36950 6010
rect 37002 5958 37014 6010
rect 37066 5958 37078 6010
rect 37130 5958 37142 6010
rect 37194 5958 37206 6010
rect 37258 5958 38824 6010
rect 1104 5936 38824 5958
rect 1104 5466 38824 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 7610 5466
rect 7662 5414 7674 5466
rect 7726 5414 7738 5466
rect 7790 5414 7802 5466
rect 7854 5414 7866 5466
rect 7918 5414 12610 5466
rect 12662 5414 12674 5466
rect 12726 5414 12738 5466
rect 12790 5414 12802 5466
rect 12854 5414 12866 5466
rect 12918 5414 17610 5466
rect 17662 5414 17674 5466
rect 17726 5414 17738 5466
rect 17790 5414 17802 5466
rect 17854 5414 17866 5466
rect 17918 5414 22610 5466
rect 22662 5414 22674 5466
rect 22726 5414 22738 5466
rect 22790 5414 22802 5466
rect 22854 5414 22866 5466
rect 22918 5414 27610 5466
rect 27662 5414 27674 5466
rect 27726 5414 27738 5466
rect 27790 5414 27802 5466
rect 27854 5414 27866 5466
rect 27918 5414 32610 5466
rect 32662 5414 32674 5466
rect 32726 5414 32738 5466
rect 32790 5414 32802 5466
rect 32854 5414 32866 5466
rect 32918 5414 37610 5466
rect 37662 5414 37674 5466
rect 37726 5414 37738 5466
rect 37790 5414 37802 5466
rect 37854 5414 37866 5466
rect 37918 5414 38824 5466
rect 1104 5392 38824 5414
rect 1104 4922 38824 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 6950 4922
rect 7002 4870 7014 4922
rect 7066 4870 7078 4922
rect 7130 4870 7142 4922
rect 7194 4870 7206 4922
rect 7258 4870 11950 4922
rect 12002 4870 12014 4922
rect 12066 4870 12078 4922
rect 12130 4870 12142 4922
rect 12194 4870 12206 4922
rect 12258 4870 16950 4922
rect 17002 4870 17014 4922
rect 17066 4870 17078 4922
rect 17130 4870 17142 4922
rect 17194 4870 17206 4922
rect 17258 4870 21950 4922
rect 22002 4870 22014 4922
rect 22066 4870 22078 4922
rect 22130 4870 22142 4922
rect 22194 4870 22206 4922
rect 22258 4870 26950 4922
rect 27002 4870 27014 4922
rect 27066 4870 27078 4922
rect 27130 4870 27142 4922
rect 27194 4870 27206 4922
rect 27258 4870 31950 4922
rect 32002 4870 32014 4922
rect 32066 4870 32078 4922
rect 32130 4870 32142 4922
rect 32194 4870 32206 4922
rect 32258 4870 36950 4922
rect 37002 4870 37014 4922
rect 37066 4870 37078 4922
rect 37130 4870 37142 4922
rect 37194 4870 37206 4922
rect 37258 4870 38824 4922
rect 1104 4848 38824 4870
rect 1104 4378 38824 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 7610 4378
rect 7662 4326 7674 4378
rect 7726 4326 7738 4378
rect 7790 4326 7802 4378
rect 7854 4326 7866 4378
rect 7918 4326 12610 4378
rect 12662 4326 12674 4378
rect 12726 4326 12738 4378
rect 12790 4326 12802 4378
rect 12854 4326 12866 4378
rect 12918 4326 17610 4378
rect 17662 4326 17674 4378
rect 17726 4326 17738 4378
rect 17790 4326 17802 4378
rect 17854 4326 17866 4378
rect 17918 4326 22610 4378
rect 22662 4326 22674 4378
rect 22726 4326 22738 4378
rect 22790 4326 22802 4378
rect 22854 4326 22866 4378
rect 22918 4326 27610 4378
rect 27662 4326 27674 4378
rect 27726 4326 27738 4378
rect 27790 4326 27802 4378
rect 27854 4326 27866 4378
rect 27918 4326 32610 4378
rect 32662 4326 32674 4378
rect 32726 4326 32738 4378
rect 32790 4326 32802 4378
rect 32854 4326 32866 4378
rect 32918 4326 37610 4378
rect 37662 4326 37674 4378
rect 37726 4326 37738 4378
rect 37790 4326 37802 4378
rect 37854 4326 37866 4378
rect 37918 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 6950 3834
rect 7002 3782 7014 3834
rect 7066 3782 7078 3834
rect 7130 3782 7142 3834
rect 7194 3782 7206 3834
rect 7258 3782 11950 3834
rect 12002 3782 12014 3834
rect 12066 3782 12078 3834
rect 12130 3782 12142 3834
rect 12194 3782 12206 3834
rect 12258 3782 16950 3834
rect 17002 3782 17014 3834
rect 17066 3782 17078 3834
rect 17130 3782 17142 3834
rect 17194 3782 17206 3834
rect 17258 3782 21950 3834
rect 22002 3782 22014 3834
rect 22066 3782 22078 3834
rect 22130 3782 22142 3834
rect 22194 3782 22206 3834
rect 22258 3782 26950 3834
rect 27002 3782 27014 3834
rect 27066 3782 27078 3834
rect 27130 3782 27142 3834
rect 27194 3782 27206 3834
rect 27258 3782 31950 3834
rect 32002 3782 32014 3834
rect 32066 3782 32078 3834
rect 32130 3782 32142 3834
rect 32194 3782 32206 3834
rect 32258 3782 36950 3834
rect 37002 3782 37014 3834
rect 37066 3782 37078 3834
rect 37130 3782 37142 3834
rect 37194 3782 37206 3834
rect 37258 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 7610 3290
rect 7662 3238 7674 3290
rect 7726 3238 7738 3290
rect 7790 3238 7802 3290
rect 7854 3238 7866 3290
rect 7918 3238 12610 3290
rect 12662 3238 12674 3290
rect 12726 3238 12738 3290
rect 12790 3238 12802 3290
rect 12854 3238 12866 3290
rect 12918 3238 17610 3290
rect 17662 3238 17674 3290
rect 17726 3238 17738 3290
rect 17790 3238 17802 3290
rect 17854 3238 17866 3290
rect 17918 3238 22610 3290
rect 22662 3238 22674 3290
rect 22726 3238 22738 3290
rect 22790 3238 22802 3290
rect 22854 3238 22866 3290
rect 22918 3238 27610 3290
rect 27662 3238 27674 3290
rect 27726 3238 27738 3290
rect 27790 3238 27802 3290
rect 27854 3238 27866 3290
rect 27918 3238 32610 3290
rect 32662 3238 32674 3290
rect 32726 3238 32738 3290
rect 32790 3238 32802 3290
rect 32854 3238 32866 3290
rect 32918 3238 37610 3290
rect 37662 3238 37674 3290
rect 37726 3238 37738 3290
rect 37790 3238 37802 3290
rect 37854 3238 37866 3290
rect 37918 3238 38824 3290
rect 1104 3216 38824 3238
rect 1104 2746 38824 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 6950 2746
rect 7002 2694 7014 2746
rect 7066 2694 7078 2746
rect 7130 2694 7142 2746
rect 7194 2694 7206 2746
rect 7258 2694 11950 2746
rect 12002 2694 12014 2746
rect 12066 2694 12078 2746
rect 12130 2694 12142 2746
rect 12194 2694 12206 2746
rect 12258 2694 16950 2746
rect 17002 2694 17014 2746
rect 17066 2694 17078 2746
rect 17130 2694 17142 2746
rect 17194 2694 17206 2746
rect 17258 2694 21950 2746
rect 22002 2694 22014 2746
rect 22066 2694 22078 2746
rect 22130 2694 22142 2746
rect 22194 2694 22206 2746
rect 22258 2694 26950 2746
rect 27002 2694 27014 2746
rect 27066 2694 27078 2746
rect 27130 2694 27142 2746
rect 27194 2694 27206 2746
rect 27258 2694 31950 2746
rect 32002 2694 32014 2746
rect 32066 2694 32078 2746
rect 32130 2694 32142 2746
rect 32194 2694 32206 2746
rect 32258 2694 36950 2746
rect 37002 2694 37014 2746
rect 37066 2694 37078 2746
rect 37130 2694 37142 2746
rect 37194 2694 37206 2746
rect 37258 2694 38824 2746
rect 1104 2672 38824 2694
rect 1104 2202 38824 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 7610 2202
rect 7662 2150 7674 2202
rect 7726 2150 7738 2202
rect 7790 2150 7802 2202
rect 7854 2150 7866 2202
rect 7918 2150 12610 2202
rect 12662 2150 12674 2202
rect 12726 2150 12738 2202
rect 12790 2150 12802 2202
rect 12854 2150 12866 2202
rect 12918 2150 17610 2202
rect 17662 2150 17674 2202
rect 17726 2150 17738 2202
rect 17790 2150 17802 2202
rect 17854 2150 17866 2202
rect 17918 2150 22610 2202
rect 22662 2150 22674 2202
rect 22726 2150 22738 2202
rect 22790 2150 22802 2202
rect 22854 2150 22866 2202
rect 22918 2150 27610 2202
rect 27662 2150 27674 2202
rect 27726 2150 27738 2202
rect 27790 2150 27802 2202
rect 27854 2150 27866 2202
rect 27918 2150 32610 2202
rect 32662 2150 32674 2202
rect 32726 2150 32738 2202
rect 32790 2150 32802 2202
rect 32854 2150 32866 2202
rect 32918 2150 37610 2202
rect 37662 2150 37674 2202
rect 37726 2150 37738 2202
rect 37790 2150 37802 2202
rect 37854 2150 37866 2202
rect 37918 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 1950 37510 2002 37562
rect 2014 37510 2066 37562
rect 2078 37510 2130 37562
rect 2142 37510 2194 37562
rect 2206 37510 2258 37562
rect 6950 37510 7002 37562
rect 7014 37510 7066 37562
rect 7078 37510 7130 37562
rect 7142 37510 7194 37562
rect 7206 37510 7258 37562
rect 11950 37510 12002 37562
rect 12014 37510 12066 37562
rect 12078 37510 12130 37562
rect 12142 37510 12194 37562
rect 12206 37510 12258 37562
rect 16950 37510 17002 37562
rect 17014 37510 17066 37562
rect 17078 37510 17130 37562
rect 17142 37510 17194 37562
rect 17206 37510 17258 37562
rect 21950 37510 22002 37562
rect 22014 37510 22066 37562
rect 22078 37510 22130 37562
rect 22142 37510 22194 37562
rect 22206 37510 22258 37562
rect 26950 37510 27002 37562
rect 27014 37510 27066 37562
rect 27078 37510 27130 37562
rect 27142 37510 27194 37562
rect 27206 37510 27258 37562
rect 31950 37510 32002 37562
rect 32014 37510 32066 37562
rect 32078 37510 32130 37562
rect 32142 37510 32194 37562
rect 32206 37510 32258 37562
rect 36950 37510 37002 37562
rect 37014 37510 37066 37562
rect 37078 37510 37130 37562
rect 37142 37510 37194 37562
rect 37206 37510 37258 37562
rect 2610 36966 2662 37018
rect 2674 36966 2726 37018
rect 2738 36966 2790 37018
rect 2802 36966 2854 37018
rect 2866 36966 2918 37018
rect 7610 36966 7662 37018
rect 7674 36966 7726 37018
rect 7738 36966 7790 37018
rect 7802 36966 7854 37018
rect 7866 36966 7918 37018
rect 12610 36966 12662 37018
rect 12674 36966 12726 37018
rect 12738 36966 12790 37018
rect 12802 36966 12854 37018
rect 12866 36966 12918 37018
rect 17610 36966 17662 37018
rect 17674 36966 17726 37018
rect 17738 36966 17790 37018
rect 17802 36966 17854 37018
rect 17866 36966 17918 37018
rect 22610 36966 22662 37018
rect 22674 36966 22726 37018
rect 22738 36966 22790 37018
rect 22802 36966 22854 37018
rect 22866 36966 22918 37018
rect 27610 36966 27662 37018
rect 27674 36966 27726 37018
rect 27738 36966 27790 37018
rect 27802 36966 27854 37018
rect 27866 36966 27918 37018
rect 32610 36966 32662 37018
rect 32674 36966 32726 37018
rect 32738 36966 32790 37018
rect 32802 36966 32854 37018
rect 32866 36966 32918 37018
rect 37610 36966 37662 37018
rect 37674 36966 37726 37018
rect 37738 36966 37790 37018
rect 37802 36966 37854 37018
rect 37866 36966 37918 37018
rect 1950 36422 2002 36474
rect 2014 36422 2066 36474
rect 2078 36422 2130 36474
rect 2142 36422 2194 36474
rect 2206 36422 2258 36474
rect 6950 36422 7002 36474
rect 7014 36422 7066 36474
rect 7078 36422 7130 36474
rect 7142 36422 7194 36474
rect 7206 36422 7258 36474
rect 11950 36422 12002 36474
rect 12014 36422 12066 36474
rect 12078 36422 12130 36474
rect 12142 36422 12194 36474
rect 12206 36422 12258 36474
rect 16950 36422 17002 36474
rect 17014 36422 17066 36474
rect 17078 36422 17130 36474
rect 17142 36422 17194 36474
rect 17206 36422 17258 36474
rect 21950 36422 22002 36474
rect 22014 36422 22066 36474
rect 22078 36422 22130 36474
rect 22142 36422 22194 36474
rect 22206 36422 22258 36474
rect 26950 36422 27002 36474
rect 27014 36422 27066 36474
rect 27078 36422 27130 36474
rect 27142 36422 27194 36474
rect 27206 36422 27258 36474
rect 31950 36422 32002 36474
rect 32014 36422 32066 36474
rect 32078 36422 32130 36474
rect 32142 36422 32194 36474
rect 32206 36422 32258 36474
rect 36950 36422 37002 36474
rect 37014 36422 37066 36474
rect 37078 36422 37130 36474
rect 37142 36422 37194 36474
rect 37206 36422 37258 36474
rect 2610 35878 2662 35930
rect 2674 35878 2726 35930
rect 2738 35878 2790 35930
rect 2802 35878 2854 35930
rect 2866 35878 2918 35930
rect 7610 35878 7662 35930
rect 7674 35878 7726 35930
rect 7738 35878 7790 35930
rect 7802 35878 7854 35930
rect 7866 35878 7918 35930
rect 12610 35878 12662 35930
rect 12674 35878 12726 35930
rect 12738 35878 12790 35930
rect 12802 35878 12854 35930
rect 12866 35878 12918 35930
rect 17610 35878 17662 35930
rect 17674 35878 17726 35930
rect 17738 35878 17790 35930
rect 17802 35878 17854 35930
rect 17866 35878 17918 35930
rect 22610 35878 22662 35930
rect 22674 35878 22726 35930
rect 22738 35878 22790 35930
rect 22802 35878 22854 35930
rect 22866 35878 22918 35930
rect 27610 35878 27662 35930
rect 27674 35878 27726 35930
rect 27738 35878 27790 35930
rect 27802 35878 27854 35930
rect 27866 35878 27918 35930
rect 32610 35878 32662 35930
rect 32674 35878 32726 35930
rect 32738 35878 32790 35930
rect 32802 35878 32854 35930
rect 32866 35878 32918 35930
rect 37610 35878 37662 35930
rect 37674 35878 37726 35930
rect 37738 35878 37790 35930
rect 37802 35878 37854 35930
rect 37866 35878 37918 35930
rect 1950 35334 2002 35386
rect 2014 35334 2066 35386
rect 2078 35334 2130 35386
rect 2142 35334 2194 35386
rect 2206 35334 2258 35386
rect 6950 35334 7002 35386
rect 7014 35334 7066 35386
rect 7078 35334 7130 35386
rect 7142 35334 7194 35386
rect 7206 35334 7258 35386
rect 11950 35334 12002 35386
rect 12014 35334 12066 35386
rect 12078 35334 12130 35386
rect 12142 35334 12194 35386
rect 12206 35334 12258 35386
rect 16950 35334 17002 35386
rect 17014 35334 17066 35386
rect 17078 35334 17130 35386
rect 17142 35334 17194 35386
rect 17206 35334 17258 35386
rect 21950 35334 22002 35386
rect 22014 35334 22066 35386
rect 22078 35334 22130 35386
rect 22142 35334 22194 35386
rect 22206 35334 22258 35386
rect 26950 35334 27002 35386
rect 27014 35334 27066 35386
rect 27078 35334 27130 35386
rect 27142 35334 27194 35386
rect 27206 35334 27258 35386
rect 31950 35334 32002 35386
rect 32014 35334 32066 35386
rect 32078 35334 32130 35386
rect 32142 35334 32194 35386
rect 32206 35334 32258 35386
rect 36950 35334 37002 35386
rect 37014 35334 37066 35386
rect 37078 35334 37130 35386
rect 37142 35334 37194 35386
rect 37206 35334 37258 35386
rect 2610 34790 2662 34842
rect 2674 34790 2726 34842
rect 2738 34790 2790 34842
rect 2802 34790 2854 34842
rect 2866 34790 2918 34842
rect 7610 34790 7662 34842
rect 7674 34790 7726 34842
rect 7738 34790 7790 34842
rect 7802 34790 7854 34842
rect 7866 34790 7918 34842
rect 12610 34790 12662 34842
rect 12674 34790 12726 34842
rect 12738 34790 12790 34842
rect 12802 34790 12854 34842
rect 12866 34790 12918 34842
rect 17610 34790 17662 34842
rect 17674 34790 17726 34842
rect 17738 34790 17790 34842
rect 17802 34790 17854 34842
rect 17866 34790 17918 34842
rect 22610 34790 22662 34842
rect 22674 34790 22726 34842
rect 22738 34790 22790 34842
rect 22802 34790 22854 34842
rect 22866 34790 22918 34842
rect 27610 34790 27662 34842
rect 27674 34790 27726 34842
rect 27738 34790 27790 34842
rect 27802 34790 27854 34842
rect 27866 34790 27918 34842
rect 32610 34790 32662 34842
rect 32674 34790 32726 34842
rect 32738 34790 32790 34842
rect 32802 34790 32854 34842
rect 32866 34790 32918 34842
rect 37610 34790 37662 34842
rect 37674 34790 37726 34842
rect 37738 34790 37790 34842
rect 37802 34790 37854 34842
rect 37866 34790 37918 34842
rect 1950 34246 2002 34298
rect 2014 34246 2066 34298
rect 2078 34246 2130 34298
rect 2142 34246 2194 34298
rect 2206 34246 2258 34298
rect 6950 34246 7002 34298
rect 7014 34246 7066 34298
rect 7078 34246 7130 34298
rect 7142 34246 7194 34298
rect 7206 34246 7258 34298
rect 11950 34246 12002 34298
rect 12014 34246 12066 34298
rect 12078 34246 12130 34298
rect 12142 34246 12194 34298
rect 12206 34246 12258 34298
rect 16950 34246 17002 34298
rect 17014 34246 17066 34298
rect 17078 34246 17130 34298
rect 17142 34246 17194 34298
rect 17206 34246 17258 34298
rect 21950 34246 22002 34298
rect 22014 34246 22066 34298
rect 22078 34246 22130 34298
rect 22142 34246 22194 34298
rect 22206 34246 22258 34298
rect 26950 34246 27002 34298
rect 27014 34246 27066 34298
rect 27078 34246 27130 34298
rect 27142 34246 27194 34298
rect 27206 34246 27258 34298
rect 31950 34246 32002 34298
rect 32014 34246 32066 34298
rect 32078 34246 32130 34298
rect 32142 34246 32194 34298
rect 32206 34246 32258 34298
rect 36950 34246 37002 34298
rect 37014 34246 37066 34298
rect 37078 34246 37130 34298
rect 37142 34246 37194 34298
rect 37206 34246 37258 34298
rect 2610 33702 2662 33754
rect 2674 33702 2726 33754
rect 2738 33702 2790 33754
rect 2802 33702 2854 33754
rect 2866 33702 2918 33754
rect 7610 33702 7662 33754
rect 7674 33702 7726 33754
rect 7738 33702 7790 33754
rect 7802 33702 7854 33754
rect 7866 33702 7918 33754
rect 12610 33702 12662 33754
rect 12674 33702 12726 33754
rect 12738 33702 12790 33754
rect 12802 33702 12854 33754
rect 12866 33702 12918 33754
rect 17610 33702 17662 33754
rect 17674 33702 17726 33754
rect 17738 33702 17790 33754
rect 17802 33702 17854 33754
rect 17866 33702 17918 33754
rect 22610 33702 22662 33754
rect 22674 33702 22726 33754
rect 22738 33702 22790 33754
rect 22802 33702 22854 33754
rect 22866 33702 22918 33754
rect 27610 33702 27662 33754
rect 27674 33702 27726 33754
rect 27738 33702 27790 33754
rect 27802 33702 27854 33754
rect 27866 33702 27918 33754
rect 32610 33702 32662 33754
rect 32674 33702 32726 33754
rect 32738 33702 32790 33754
rect 32802 33702 32854 33754
rect 32866 33702 32918 33754
rect 37610 33702 37662 33754
rect 37674 33702 37726 33754
rect 37738 33702 37790 33754
rect 37802 33702 37854 33754
rect 37866 33702 37918 33754
rect 1950 33158 2002 33210
rect 2014 33158 2066 33210
rect 2078 33158 2130 33210
rect 2142 33158 2194 33210
rect 2206 33158 2258 33210
rect 6950 33158 7002 33210
rect 7014 33158 7066 33210
rect 7078 33158 7130 33210
rect 7142 33158 7194 33210
rect 7206 33158 7258 33210
rect 11950 33158 12002 33210
rect 12014 33158 12066 33210
rect 12078 33158 12130 33210
rect 12142 33158 12194 33210
rect 12206 33158 12258 33210
rect 16950 33158 17002 33210
rect 17014 33158 17066 33210
rect 17078 33158 17130 33210
rect 17142 33158 17194 33210
rect 17206 33158 17258 33210
rect 21950 33158 22002 33210
rect 22014 33158 22066 33210
rect 22078 33158 22130 33210
rect 22142 33158 22194 33210
rect 22206 33158 22258 33210
rect 26950 33158 27002 33210
rect 27014 33158 27066 33210
rect 27078 33158 27130 33210
rect 27142 33158 27194 33210
rect 27206 33158 27258 33210
rect 31950 33158 32002 33210
rect 32014 33158 32066 33210
rect 32078 33158 32130 33210
rect 32142 33158 32194 33210
rect 32206 33158 32258 33210
rect 36950 33158 37002 33210
rect 37014 33158 37066 33210
rect 37078 33158 37130 33210
rect 37142 33158 37194 33210
rect 37206 33158 37258 33210
rect 2610 32614 2662 32666
rect 2674 32614 2726 32666
rect 2738 32614 2790 32666
rect 2802 32614 2854 32666
rect 2866 32614 2918 32666
rect 7610 32614 7662 32666
rect 7674 32614 7726 32666
rect 7738 32614 7790 32666
rect 7802 32614 7854 32666
rect 7866 32614 7918 32666
rect 12610 32614 12662 32666
rect 12674 32614 12726 32666
rect 12738 32614 12790 32666
rect 12802 32614 12854 32666
rect 12866 32614 12918 32666
rect 17610 32614 17662 32666
rect 17674 32614 17726 32666
rect 17738 32614 17790 32666
rect 17802 32614 17854 32666
rect 17866 32614 17918 32666
rect 22610 32614 22662 32666
rect 22674 32614 22726 32666
rect 22738 32614 22790 32666
rect 22802 32614 22854 32666
rect 22866 32614 22918 32666
rect 27610 32614 27662 32666
rect 27674 32614 27726 32666
rect 27738 32614 27790 32666
rect 27802 32614 27854 32666
rect 27866 32614 27918 32666
rect 32610 32614 32662 32666
rect 32674 32614 32726 32666
rect 32738 32614 32790 32666
rect 32802 32614 32854 32666
rect 32866 32614 32918 32666
rect 37610 32614 37662 32666
rect 37674 32614 37726 32666
rect 37738 32614 37790 32666
rect 37802 32614 37854 32666
rect 37866 32614 37918 32666
rect 1950 32070 2002 32122
rect 2014 32070 2066 32122
rect 2078 32070 2130 32122
rect 2142 32070 2194 32122
rect 2206 32070 2258 32122
rect 6950 32070 7002 32122
rect 7014 32070 7066 32122
rect 7078 32070 7130 32122
rect 7142 32070 7194 32122
rect 7206 32070 7258 32122
rect 11950 32070 12002 32122
rect 12014 32070 12066 32122
rect 12078 32070 12130 32122
rect 12142 32070 12194 32122
rect 12206 32070 12258 32122
rect 16950 32070 17002 32122
rect 17014 32070 17066 32122
rect 17078 32070 17130 32122
rect 17142 32070 17194 32122
rect 17206 32070 17258 32122
rect 21950 32070 22002 32122
rect 22014 32070 22066 32122
rect 22078 32070 22130 32122
rect 22142 32070 22194 32122
rect 22206 32070 22258 32122
rect 26950 32070 27002 32122
rect 27014 32070 27066 32122
rect 27078 32070 27130 32122
rect 27142 32070 27194 32122
rect 27206 32070 27258 32122
rect 31950 32070 32002 32122
rect 32014 32070 32066 32122
rect 32078 32070 32130 32122
rect 32142 32070 32194 32122
rect 32206 32070 32258 32122
rect 36950 32070 37002 32122
rect 37014 32070 37066 32122
rect 37078 32070 37130 32122
rect 37142 32070 37194 32122
rect 37206 32070 37258 32122
rect 2610 31526 2662 31578
rect 2674 31526 2726 31578
rect 2738 31526 2790 31578
rect 2802 31526 2854 31578
rect 2866 31526 2918 31578
rect 7610 31526 7662 31578
rect 7674 31526 7726 31578
rect 7738 31526 7790 31578
rect 7802 31526 7854 31578
rect 7866 31526 7918 31578
rect 12610 31526 12662 31578
rect 12674 31526 12726 31578
rect 12738 31526 12790 31578
rect 12802 31526 12854 31578
rect 12866 31526 12918 31578
rect 17610 31526 17662 31578
rect 17674 31526 17726 31578
rect 17738 31526 17790 31578
rect 17802 31526 17854 31578
rect 17866 31526 17918 31578
rect 22610 31526 22662 31578
rect 22674 31526 22726 31578
rect 22738 31526 22790 31578
rect 22802 31526 22854 31578
rect 22866 31526 22918 31578
rect 27610 31526 27662 31578
rect 27674 31526 27726 31578
rect 27738 31526 27790 31578
rect 27802 31526 27854 31578
rect 27866 31526 27918 31578
rect 32610 31526 32662 31578
rect 32674 31526 32726 31578
rect 32738 31526 32790 31578
rect 32802 31526 32854 31578
rect 32866 31526 32918 31578
rect 37610 31526 37662 31578
rect 37674 31526 37726 31578
rect 37738 31526 37790 31578
rect 37802 31526 37854 31578
rect 37866 31526 37918 31578
rect 1950 30982 2002 31034
rect 2014 30982 2066 31034
rect 2078 30982 2130 31034
rect 2142 30982 2194 31034
rect 2206 30982 2258 31034
rect 6950 30982 7002 31034
rect 7014 30982 7066 31034
rect 7078 30982 7130 31034
rect 7142 30982 7194 31034
rect 7206 30982 7258 31034
rect 11950 30982 12002 31034
rect 12014 30982 12066 31034
rect 12078 30982 12130 31034
rect 12142 30982 12194 31034
rect 12206 30982 12258 31034
rect 16950 30982 17002 31034
rect 17014 30982 17066 31034
rect 17078 30982 17130 31034
rect 17142 30982 17194 31034
rect 17206 30982 17258 31034
rect 21950 30982 22002 31034
rect 22014 30982 22066 31034
rect 22078 30982 22130 31034
rect 22142 30982 22194 31034
rect 22206 30982 22258 31034
rect 26950 30982 27002 31034
rect 27014 30982 27066 31034
rect 27078 30982 27130 31034
rect 27142 30982 27194 31034
rect 27206 30982 27258 31034
rect 31950 30982 32002 31034
rect 32014 30982 32066 31034
rect 32078 30982 32130 31034
rect 32142 30982 32194 31034
rect 32206 30982 32258 31034
rect 36950 30982 37002 31034
rect 37014 30982 37066 31034
rect 37078 30982 37130 31034
rect 37142 30982 37194 31034
rect 37206 30982 37258 31034
rect 2610 30438 2662 30490
rect 2674 30438 2726 30490
rect 2738 30438 2790 30490
rect 2802 30438 2854 30490
rect 2866 30438 2918 30490
rect 7610 30438 7662 30490
rect 7674 30438 7726 30490
rect 7738 30438 7790 30490
rect 7802 30438 7854 30490
rect 7866 30438 7918 30490
rect 12610 30438 12662 30490
rect 12674 30438 12726 30490
rect 12738 30438 12790 30490
rect 12802 30438 12854 30490
rect 12866 30438 12918 30490
rect 17610 30438 17662 30490
rect 17674 30438 17726 30490
rect 17738 30438 17790 30490
rect 17802 30438 17854 30490
rect 17866 30438 17918 30490
rect 22610 30438 22662 30490
rect 22674 30438 22726 30490
rect 22738 30438 22790 30490
rect 22802 30438 22854 30490
rect 22866 30438 22918 30490
rect 27610 30438 27662 30490
rect 27674 30438 27726 30490
rect 27738 30438 27790 30490
rect 27802 30438 27854 30490
rect 27866 30438 27918 30490
rect 32610 30438 32662 30490
rect 32674 30438 32726 30490
rect 32738 30438 32790 30490
rect 32802 30438 32854 30490
rect 32866 30438 32918 30490
rect 37610 30438 37662 30490
rect 37674 30438 37726 30490
rect 37738 30438 37790 30490
rect 37802 30438 37854 30490
rect 37866 30438 37918 30490
rect 1950 29894 2002 29946
rect 2014 29894 2066 29946
rect 2078 29894 2130 29946
rect 2142 29894 2194 29946
rect 2206 29894 2258 29946
rect 6950 29894 7002 29946
rect 7014 29894 7066 29946
rect 7078 29894 7130 29946
rect 7142 29894 7194 29946
rect 7206 29894 7258 29946
rect 11950 29894 12002 29946
rect 12014 29894 12066 29946
rect 12078 29894 12130 29946
rect 12142 29894 12194 29946
rect 12206 29894 12258 29946
rect 16950 29894 17002 29946
rect 17014 29894 17066 29946
rect 17078 29894 17130 29946
rect 17142 29894 17194 29946
rect 17206 29894 17258 29946
rect 21950 29894 22002 29946
rect 22014 29894 22066 29946
rect 22078 29894 22130 29946
rect 22142 29894 22194 29946
rect 22206 29894 22258 29946
rect 26950 29894 27002 29946
rect 27014 29894 27066 29946
rect 27078 29894 27130 29946
rect 27142 29894 27194 29946
rect 27206 29894 27258 29946
rect 31950 29894 32002 29946
rect 32014 29894 32066 29946
rect 32078 29894 32130 29946
rect 32142 29894 32194 29946
rect 32206 29894 32258 29946
rect 36950 29894 37002 29946
rect 37014 29894 37066 29946
rect 37078 29894 37130 29946
rect 37142 29894 37194 29946
rect 37206 29894 37258 29946
rect 2610 29350 2662 29402
rect 2674 29350 2726 29402
rect 2738 29350 2790 29402
rect 2802 29350 2854 29402
rect 2866 29350 2918 29402
rect 7610 29350 7662 29402
rect 7674 29350 7726 29402
rect 7738 29350 7790 29402
rect 7802 29350 7854 29402
rect 7866 29350 7918 29402
rect 12610 29350 12662 29402
rect 12674 29350 12726 29402
rect 12738 29350 12790 29402
rect 12802 29350 12854 29402
rect 12866 29350 12918 29402
rect 17610 29350 17662 29402
rect 17674 29350 17726 29402
rect 17738 29350 17790 29402
rect 17802 29350 17854 29402
rect 17866 29350 17918 29402
rect 22610 29350 22662 29402
rect 22674 29350 22726 29402
rect 22738 29350 22790 29402
rect 22802 29350 22854 29402
rect 22866 29350 22918 29402
rect 27610 29350 27662 29402
rect 27674 29350 27726 29402
rect 27738 29350 27790 29402
rect 27802 29350 27854 29402
rect 27866 29350 27918 29402
rect 32610 29350 32662 29402
rect 32674 29350 32726 29402
rect 32738 29350 32790 29402
rect 32802 29350 32854 29402
rect 32866 29350 32918 29402
rect 37610 29350 37662 29402
rect 37674 29350 37726 29402
rect 37738 29350 37790 29402
rect 37802 29350 37854 29402
rect 37866 29350 37918 29402
rect 1950 28806 2002 28858
rect 2014 28806 2066 28858
rect 2078 28806 2130 28858
rect 2142 28806 2194 28858
rect 2206 28806 2258 28858
rect 6950 28806 7002 28858
rect 7014 28806 7066 28858
rect 7078 28806 7130 28858
rect 7142 28806 7194 28858
rect 7206 28806 7258 28858
rect 11950 28806 12002 28858
rect 12014 28806 12066 28858
rect 12078 28806 12130 28858
rect 12142 28806 12194 28858
rect 12206 28806 12258 28858
rect 16950 28806 17002 28858
rect 17014 28806 17066 28858
rect 17078 28806 17130 28858
rect 17142 28806 17194 28858
rect 17206 28806 17258 28858
rect 21950 28806 22002 28858
rect 22014 28806 22066 28858
rect 22078 28806 22130 28858
rect 22142 28806 22194 28858
rect 22206 28806 22258 28858
rect 26950 28806 27002 28858
rect 27014 28806 27066 28858
rect 27078 28806 27130 28858
rect 27142 28806 27194 28858
rect 27206 28806 27258 28858
rect 31950 28806 32002 28858
rect 32014 28806 32066 28858
rect 32078 28806 32130 28858
rect 32142 28806 32194 28858
rect 32206 28806 32258 28858
rect 36950 28806 37002 28858
rect 37014 28806 37066 28858
rect 37078 28806 37130 28858
rect 37142 28806 37194 28858
rect 37206 28806 37258 28858
rect 2610 28262 2662 28314
rect 2674 28262 2726 28314
rect 2738 28262 2790 28314
rect 2802 28262 2854 28314
rect 2866 28262 2918 28314
rect 7610 28262 7662 28314
rect 7674 28262 7726 28314
rect 7738 28262 7790 28314
rect 7802 28262 7854 28314
rect 7866 28262 7918 28314
rect 12610 28262 12662 28314
rect 12674 28262 12726 28314
rect 12738 28262 12790 28314
rect 12802 28262 12854 28314
rect 12866 28262 12918 28314
rect 17610 28262 17662 28314
rect 17674 28262 17726 28314
rect 17738 28262 17790 28314
rect 17802 28262 17854 28314
rect 17866 28262 17918 28314
rect 22610 28262 22662 28314
rect 22674 28262 22726 28314
rect 22738 28262 22790 28314
rect 22802 28262 22854 28314
rect 22866 28262 22918 28314
rect 27610 28262 27662 28314
rect 27674 28262 27726 28314
rect 27738 28262 27790 28314
rect 27802 28262 27854 28314
rect 27866 28262 27918 28314
rect 32610 28262 32662 28314
rect 32674 28262 32726 28314
rect 32738 28262 32790 28314
rect 32802 28262 32854 28314
rect 32866 28262 32918 28314
rect 37610 28262 37662 28314
rect 37674 28262 37726 28314
rect 37738 28262 37790 28314
rect 37802 28262 37854 28314
rect 37866 28262 37918 28314
rect 1950 27718 2002 27770
rect 2014 27718 2066 27770
rect 2078 27718 2130 27770
rect 2142 27718 2194 27770
rect 2206 27718 2258 27770
rect 6950 27718 7002 27770
rect 7014 27718 7066 27770
rect 7078 27718 7130 27770
rect 7142 27718 7194 27770
rect 7206 27718 7258 27770
rect 11950 27718 12002 27770
rect 12014 27718 12066 27770
rect 12078 27718 12130 27770
rect 12142 27718 12194 27770
rect 12206 27718 12258 27770
rect 16950 27718 17002 27770
rect 17014 27718 17066 27770
rect 17078 27718 17130 27770
rect 17142 27718 17194 27770
rect 17206 27718 17258 27770
rect 21950 27718 22002 27770
rect 22014 27718 22066 27770
rect 22078 27718 22130 27770
rect 22142 27718 22194 27770
rect 22206 27718 22258 27770
rect 26950 27718 27002 27770
rect 27014 27718 27066 27770
rect 27078 27718 27130 27770
rect 27142 27718 27194 27770
rect 27206 27718 27258 27770
rect 31950 27718 32002 27770
rect 32014 27718 32066 27770
rect 32078 27718 32130 27770
rect 32142 27718 32194 27770
rect 32206 27718 32258 27770
rect 36950 27718 37002 27770
rect 37014 27718 37066 27770
rect 37078 27718 37130 27770
rect 37142 27718 37194 27770
rect 37206 27718 37258 27770
rect 2610 27174 2662 27226
rect 2674 27174 2726 27226
rect 2738 27174 2790 27226
rect 2802 27174 2854 27226
rect 2866 27174 2918 27226
rect 7610 27174 7662 27226
rect 7674 27174 7726 27226
rect 7738 27174 7790 27226
rect 7802 27174 7854 27226
rect 7866 27174 7918 27226
rect 12610 27174 12662 27226
rect 12674 27174 12726 27226
rect 12738 27174 12790 27226
rect 12802 27174 12854 27226
rect 12866 27174 12918 27226
rect 17610 27174 17662 27226
rect 17674 27174 17726 27226
rect 17738 27174 17790 27226
rect 17802 27174 17854 27226
rect 17866 27174 17918 27226
rect 22610 27174 22662 27226
rect 22674 27174 22726 27226
rect 22738 27174 22790 27226
rect 22802 27174 22854 27226
rect 22866 27174 22918 27226
rect 27610 27174 27662 27226
rect 27674 27174 27726 27226
rect 27738 27174 27790 27226
rect 27802 27174 27854 27226
rect 27866 27174 27918 27226
rect 32610 27174 32662 27226
rect 32674 27174 32726 27226
rect 32738 27174 32790 27226
rect 32802 27174 32854 27226
rect 32866 27174 32918 27226
rect 37610 27174 37662 27226
rect 37674 27174 37726 27226
rect 37738 27174 37790 27226
rect 37802 27174 37854 27226
rect 37866 27174 37918 27226
rect 1950 26630 2002 26682
rect 2014 26630 2066 26682
rect 2078 26630 2130 26682
rect 2142 26630 2194 26682
rect 2206 26630 2258 26682
rect 6950 26630 7002 26682
rect 7014 26630 7066 26682
rect 7078 26630 7130 26682
rect 7142 26630 7194 26682
rect 7206 26630 7258 26682
rect 11950 26630 12002 26682
rect 12014 26630 12066 26682
rect 12078 26630 12130 26682
rect 12142 26630 12194 26682
rect 12206 26630 12258 26682
rect 16950 26630 17002 26682
rect 17014 26630 17066 26682
rect 17078 26630 17130 26682
rect 17142 26630 17194 26682
rect 17206 26630 17258 26682
rect 21950 26630 22002 26682
rect 22014 26630 22066 26682
rect 22078 26630 22130 26682
rect 22142 26630 22194 26682
rect 22206 26630 22258 26682
rect 26950 26630 27002 26682
rect 27014 26630 27066 26682
rect 27078 26630 27130 26682
rect 27142 26630 27194 26682
rect 27206 26630 27258 26682
rect 31950 26630 32002 26682
rect 32014 26630 32066 26682
rect 32078 26630 32130 26682
rect 32142 26630 32194 26682
rect 32206 26630 32258 26682
rect 36950 26630 37002 26682
rect 37014 26630 37066 26682
rect 37078 26630 37130 26682
rect 37142 26630 37194 26682
rect 37206 26630 37258 26682
rect 2610 26086 2662 26138
rect 2674 26086 2726 26138
rect 2738 26086 2790 26138
rect 2802 26086 2854 26138
rect 2866 26086 2918 26138
rect 7610 26086 7662 26138
rect 7674 26086 7726 26138
rect 7738 26086 7790 26138
rect 7802 26086 7854 26138
rect 7866 26086 7918 26138
rect 12610 26086 12662 26138
rect 12674 26086 12726 26138
rect 12738 26086 12790 26138
rect 12802 26086 12854 26138
rect 12866 26086 12918 26138
rect 17610 26086 17662 26138
rect 17674 26086 17726 26138
rect 17738 26086 17790 26138
rect 17802 26086 17854 26138
rect 17866 26086 17918 26138
rect 22610 26086 22662 26138
rect 22674 26086 22726 26138
rect 22738 26086 22790 26138
rect 22802 26086 22854 26138
rect 22866 26086 22918 26138
rect 27610 26086 27662 26138
rect 27674 26086 27726 26138
rect 27738 26086 27790 26138
rect 27802 26086 27854 26138
rect 27866 26086 27918 26138
rect 32610 26086 32662 26138
rect 32674 26086 32726 26138
rect 32738 26086 32790 26138
rect 32802 26086 32854 26138
rect 32866 26086 32918 26138
rect 37610 26086 37662 26138
rect 37674 26086 37726 26138
rect 37738 26086 37790 26138
rect 37802 26086 37854 26138
rect 37866 26086 37918 26138
rect 1950 25542 2002 25594
rect 2014 25542 2066 25594
rect 2078 25542 2130 25594
rect 2142 25542 2194 25594
rect 2206 25542 2258 25594
rect 6950 25542 7002 25594
rect 7014 25542 7066 25594
rect 7078 25542 7130 25594
rect 7142 25542 7194 25594
rect 7206 25542 7258 25594
rect 11950 25542 12002 25594
rect 12014 25542 12066 25594
rect 12078 25542 12130 25594
rect 12142 25542 12194 25594
rect 12206 25542 12258 25594
rect 16950 25542 17002 25594
rect 17014 25542 17066 25594
rect 17078 25542 17130 25594
rect 17142 25542 17194 25594
rect 17206 25542 17258 25594
rect 21950 25542 22002 25594
rect 22014 25542 22066 25594
rect 22078 25542 22130 25594
rect 22142 25542 22194 25594
rect 22206 25542 22258 25594
rect 26950 25542 27002 25594
rect 27014 25542 27066 25594
rect 27078 25542 27130 25594
rect 27142 25542 27194 25594
rect 27206 25542 27258 25594
rect 31950 25542 32002 25594
rect 32014 25542 32066 25594
rect 32078 25542 32130 25594
rect 32142 25542 32194 25594
rect 32206 25542 32258 25594
rect 36950 25542 37002 25594
rect 37014 25542 37066 25594
rect 37078 25542 37130 25594
rect 37142 25542 37194 25594
rect 37206 25542 37258 25594
rect 2610 24998 2662 25050
rect 2674 24998 2726 25050
rect 2738 24998 2790 25050
rect 2802 24998 2854 25050
rect 2866 24998 2918 25050
rect 7610 24998 7662 25050
rect 7674 24998 7726 25050
rect 7738 24998 7790 25050
rect 7802 24998 7854 25050
rect 7866 24998 7918 25050
rect 12610 24998 12662 25050
rect 12674 24998 12726 25050
rect 12738 24998 12790 25050
rect 12802 24998 12854 25050
rect 12866 24998 12918 25050
rect 17610 24998 17662 25050
rect 17674 24998 17726 25050
rect 17738 24998 17790 25050
rect 17802 24998 17854 25050
rect 17866 24998 17918 25050
rect 22610 24998 22662 25050
rect 22674 24998 22726 25050
rect 22738 24998 22790 25050
rect 22802 24998 22854 25050
rect 22866 24998 22918 25050
rect 27610 24998 27662 25050
rect 27674 24998 27726 25050
rect 27738 24998 27790 25050
rect 27802 24998 27854 25050
rect 27866 24998 27918 25050
rect 32610 24998 32662 25050
rect 32674 24998 32726 25050
rect 32738 24998 32790 25050
rect 32802 24998 32854 25050
rect 32866 24998 32918 25050
rect 37610 24998 37662 25050
rect 37674 24998 37726 25050
rect 37738 24998 37790 25050
rect 37802 24998 37854 25050
rect 37866 24998 37918 25050
rect 1950 24454 2002 24506
rect 2014 24454 2066 24506
rect 2078 24454 2130 24506
rect 2142 24454 2194 24506
rect 2206 24454 2258 24506
rect 6950 24454 7002 24506
rect 7014 24454 7066 24506
rect 7078 24454 7130 24506
rect 7142 24454 7194 24506
rect 7206 24454 7258 24506
rect 11950 24454 12002 24506
rect 12014 24454 12066 24506
rect 12078 24454 12130 24506
rect 12142 24454 12194 24506
rect 12206 24454 12258 24506
rect 16950 24454 17002 24506
rect 17014 24454 17066 24506
rect 17078 24454 17130 24506
rect 17142 24454 17194 24506
rect 17206 24454 17258 24506
rect 21950 24454 22002 24506
rect 22014 24454 22066 24506
rect 22078 24454 22130 24506
rect 22142 24454 22194 24506
rect 22206 24454 22258 24506
rect 26950 24454 27002 24506
rect 27014 24454 27066 24506
rect 27078 24454 27130 24506
rect 27142 24454 27194 24506
rect 27206 24454 27258 24506
rect 31950 24454 32002 24506
rect 32014 24454 32066 24506
rect 32078 24454 32130 24506
rect 32142 24454 32194 24506
rect 32206 24454 32258 24506
rect 36950 24454 37002 24506
rect 37014 24454 37066 24506
rect 37078 24454 37130 24506
rect 37142 24454 37194 24506
rect 37206 24454 37258 24506
rect 2610 23910 2662 23962
rect 2674 23910 2726 23962
rect 2738 23910 2790 23962
rect 2802 23910 2854 23962
rect 2866 23910 2918 23962
rect 7610 23910 7662 23962
rect 7674 23910 7726 23962
rect 7738 23910 7790 23962
rect 7802 23910 7854 23962
rect 7866 23910 7918 23962
rect 12610 23910 12662 23962
rect 12674 23910 12726 23962
rect 12738 23910 12790 23962
rect 12802 23910 12854 23962
rect 12866 23910 12918 23962
rect 17610 23910 17662 23962
rect 17674 23910 17726 23962
rect 17738 23910 17790 23962
rect 17802 23910 17854 23962
rect 17866 23910 17918 23962
rect 22610 23910 22662 23962
rect 22674 23910 22726 23962
rect 22738 23910 22790 23962
rect 22802 23910 22854 23962
rect 22866 23910 22918 23962
rect 27610 23910 27662 23962
rect 27674 23910 27726 23962
rect 27738 23910 27790 23962
rect 27802 23910 27854 23962
rect 27866 23910 27918 23962
rect 32610 23910 32662 23962
rect 32674 23910 32726 23962
rect 32738 23910 32790 23962
rect 32802 23910 32854 23962
rect 32866 23910 32918 23962
rect 37610 23910 37662 23962
rect 37674 23910 37726 23962
rect 37738 23910 37790 23962
rect 37802 23910 37854 23962
rect 37866 23910 37918 23962
rect 1950 23366 2002 23418
rect 2014 23366 2066 23418
rect 2078 23366 2130 23418
rect 2142 23366 2194 23418
rect 2206 23366 2258 23418
rect 6950 23366 7002 23418
rect 7014 23366 7066 23418
rect 7078 23366 7130 23418
rect 7142 23366 7194 23418
rect 7206 23366 7258 23418
rect 11950 23366 12002 23418
rect 12014 23366 12066 23418
rect 12078 23366 12130 23418
rect 12142 23366 12194 23418
rect 12206 23366 12258 23418
rect 16950 23366 17002 23418
rect 17014 23366 17066 23418
rect 17078 23366 17130 23418
rect 17142 23366 17194 23418
rect 17206 23366 17258 23418
rect 21950 23366 22002 23418
rect 22014 23366 22066 23418
rect 22078 23366 22130 23418
rect 22142 23366 22194 23418
rect 22206 23366 22258 23418
rect 26950 23366 27002 23418
rect 27014 23366 27066 23418
rect 27078 23366 27130 23418
rect 27142 23366 27194 23418
rect 27206 23366 27258 23418
rect 31950 23366 32002 23418
rect 32014 23366 32066 23418
rect 32078 23366 32130 23418
rect 32142 23366 32194 23418
rect 32206 23366 32258 23418
rect 36950 23366 37002 23418
rect 37014 23366 37066 23418
rect 37078 23366 37130 23418
rect 37142 23366 37194 23418
rect 37206 23366 37258 23418
rect 2610 22822 2662 22874
rect 2674 22822 2726 22874
rect 2738 22822 2790 22874
rect 2802 22822 2854 22874
rect 2866 22822 2918 22874
rect 7610 22822 7662 22874
rect 7674 22822 7726 22874
rect 7738 22822 7790 22874
rect 7802 22822 7854 22874
rect 7866 22822 7918 22874
rect 12610 22822 12662 22874
rect 12674 22822 12726 22874
rect 12738 22822 12790 22874
rect 12802 22822 12854 22874
rect 12866 22822 12918 22874
rect 17610 22822 17662 22874
rect 17674 22822 17726 22874
rect 17738 22822 17790 22874
rect 17802 22822 17854 22874
rect 17866 22822 17918 22874
rect 22610 22822 22662 22874
rect 22674 22822 22726 22874
rect 22738 22822 22790 22874
rect 22802 22822 22854 22874
rect 22866 22822 22918 22874
rect 27610 22822 27662 22874
rect 27674 22822 27726 22874
rect 27738 22822 27790 22874
rect 27802 22822 27854 22874
rect 27866 22822 27918 22874
rect 32610 22822 32662 22874
rect 32674 22822 32726 22874
rect 32738 22822 32790 22874
rect 32802 22822 32854 22874
rect 32866 22822 32918 22874
rect 37610 22822 37662 22874
rect 37674 22822 37726 22874
rect 37738 22822 37790 22874
rect 37802 22822 37854 22874
rect 37866 22822 37918 22874
rect 1950 22278 2002 22330
rect 2014 22278 2066 22330
rect 2078 22278 2130 22330
rect 2142 22278 2194 22330
rect 2206 22278 2258 22330
rect 6950 22278 7002 22330
rect 7014 22278 7066 22330
rect 7078 22278 7130 22330
rect 7142 22278 7194 22330
rect 7206 22278 7258 22330
rect 11950 22278 12002 22330
rect 12014 22278 12066 22330
rect 12078 22278 12130 22330
rect 12142 22278 12194 22330
rect 12206 22278 12258 22330
rect 16950 22278 17002 22330
rect 17014 22278 17066 22330
rect 17078 22278 17130 22330
rect 17142 22278 17194 22330
rect 17206 22278 17258 22330
rect 21950 22278 22002 22330
rect 22014 22278 22066 22330
rect 22078 22278 22130 22330
rect 22142 22278 22194 22330
rect 22206 22278 22258 22330
rect 26950 22278 27002 22330
rect 27014 22278 27066 22330
rect 27078 22278 27130 22330
rect 27142 22278 27194 22330
rect 27206 22278 27258 22330
rect 31950 22278 32002 22330
rect 32014 22278 32066 22330
rect 32078 22278 32130 22330
rect 32142 22278 32194 22330
rect 32206 22278 32258 22330
rect 36950 22278 37002 22330
rect 37014 22278 37066 22330
rect 37078 22278 37130 22330
rect 37142 22278 37194 22330
rect 37206 22278 37258 22330
rect 37280 21972 37332 22024
rect 38476 21879 38528 21888
rect 38476 21845 38485 21879
rect 38485 21845 38519 21879
rect 38519 21845 38528 21879
rect 38476 21836 38528 21845
rect 2610 21734 2662 21786
rect 2674 21734 2726 21786
rect 2738 21734 2790 21786
rect 2802 21734 2854 21786
rect 2866 21734 2918 21786
rect 7610 21734 7662 21786
rect 7674 21734 7726 21786
rect 7738 21734 7790 21786
rect 7802 21734 7854 21786
rect 7866 21734 7918 21786
rect 12610 21734 12662 21786
rect 12674 21734 12726 21786
rect 12738 21734 12790 21786
rect 12802 21734 12854 21786
rect 12866 21734 12918 21786
rect 17610 21734 17662 21786
rect 17674 21734 17726 21786
rect 17738 21734 17790 21786
rect 17802 21734 17854 21786
rect 17866 21734 17918 21786
rect 22610 21734 22662 21786
rect 22674 21734 22726 21786
rect 22738 21734 22790 21786
rect 22802 21734 22854 21786
rect 22866 21734 22918 21786
rect 27610 21734 27662 21786
rect 27674 21734 27726 21786
rect 27738 21734 27790 21786
rect 27802 21734 27854 21786
rect 27866 21734 27918 21786
rect 32610 21734 32662 21786
rect 32674 21734 32726 21786
rect 32738 21734 32790 21786
rect 32802 21734 32854 21786
rect 32866 21734 32918 21786
rect 37610 21734 37662 21786
rect 37674 21734 37726 21786
rect 37738 21734 37790 21786
rect 37802 21734 37854 21786
rect 37866 21734 37918 21786
rect 940 21496 992 21548
rect 20444 21539 20496 21548
rect 20444 21505 20453 21539
rect 20453 21505 20487 21539
rect 20487 21505 20496 21539
rect 20444 21496 20496 21505
rect 38292 21539 38344 21548
rect 38292 21505 38301 21539
rect 38301 21505 38335 21539
rect 38335 21505 38344 21539
rect 38292 21496 38344 21505
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 19800 21292 19852 21344
rect 38476 21335 38528 21344
rect 38476 21301 38485 21335
rect 38485 21301 38519 21335
rect 38519 21301 38528 21335
rect 38476 21292 38528 21301
rect 1950 21190 2002 21242
rect 2014 21190 2066 21242
rect 2078 21190 2130 21242
rect 2142 21190 2194 21242
rect 2206 21190 2258 21242
rect 6950 21190 7002 21242
rect 7014 21190 7066 21242
rect 7078 21190 7130 21242
rect 7142 21190 7194 21242
rect 7206 21190 7258 21242
rect 11950 21190 12002 21242
rect 12014 21190 12066 21242
rect 12078 21190 12130 21242
rect 12142 21190 12194 21242
rect 12206 21190 12258 21242
rect 16950 21190 17002 21242
rect 17014 21190 17066 21242
rect 17078 21190 17130 21242
rect 17142 21190 17194 21242
rect 17206 21190 17258 21242
rect 21950 21190 22002 21242
rect 22014 21190 22066 21242
rect 22078 21190 22130 21242
rect 22142 21190 22194 21242
rect 22206 21190 22258 21242
rect 26950 21190 27002 21242
rect 27014 21190 27066 21242
rect 27078 21190 27130 21242
rect 27142 21190 27194 21242
rect 27206 21190 27258 21242
rect 31950 21190 32002 21242
rect 32014 21190 32066 21242
rect 32078 21190 32130 21242
rect 32142 21190 32194 21242
rect 32206 21190 32258 21242
rect 36950 21190 37002 21242
rect 37014 21190 37066 21242
rect 37078 21190 37130 21242
rect 37142 21190 37194 21242
rect 37206 21190 37258 21242
rect 1584 21088 1636 21140
rect 15292 21088 15344 21140
rect 19800 20995 19852 21004
rect 19800 20961 19809 20995
rect 19809 20961 19843 20995
rect 19843 20961 19852 20995
rect 19800 20952 19852 20961
rect 15200 20884 15252 20936
rect 19892 20884 19944 20936
rect 34520 20884 34572 20936
rect 19708 20816 19760 20868
rect 20260 20859 20312 20868
rect 20260 20825 20269 20859
rect 20269 20825 20303 20859
rect 20303 20825 20312 20859
rect 20260 20816 20312 20825
rect 1400 20791 1452 20800
rect 1400 20757 1409 20791
rect 1409 20757 1443 20791
rect 1443 20757 1452 20791
rect 1400 20748 1452 20757
rect 20168 20748 20220 20800
rect 2610 20646 2662 20698
rect 2674 20646 2726 20698
rect 2738 20646 2790 20698
rect 2802 20646 2854 20698
rect 2866 20646 2918 20698
rect 7610 20646 7662 20698
rect 7674 20646 7726 20698
rect 7738 20646 7790 20698
rect 7802 20646 7854 20698
rect 7866 20646 7918 20698
rect 12610 20646 12662 20698
rect 12674 20646 12726 20698
rect 12738 20646 12790 20698
rect 12802 20646 12854 20698
rect 12866 20646 12918 20698
rect 17610 20646 17662 20698
rect 17674 20646 17726 20698
rect 17738 20646 17790 20698
rect 17802 20646 17854 20698
rect 17866 20646 17918 20698
rect 22610 20646 22662 20698
rect 22674 20646 22726 20698
rect 22738 20646 22790 20698
rect 22802 20646 22854 20698
rect 22866 20646 22918 20698
rect 27610 20646 27662 20698
rect 27674 20646 27726 20698
rect 27738 20646 27790 20698
rect 27802 20646 27854 20698
rect 27866 20646 27918 20698
rect 32610 20646 32662 20698
rect 32674 20646 32726 20698
rect 32738 20646 32790 20698
rect 32802 20646 32854 20698
rect 32866 20646 32918 20698
rect 37610 20646 37662 20698
rect 37674 20646 37726 20698
rect 37738 20646 37790 20698
rect 37802 20646 37854 20698
rect 37866 20646 37918 20698
rect 39028 20680 39080 20732
rect 15200 20544 15252 20596
rect 19800 20544 19852 20596
rect 20260 20544 20312 20596
rect 19432 20451 19484 20460
rect 19432 20417 19441 20451
rect 19441 20417 19475 20451
rect 19475 20417 19484 20451
rect 19432 20408 19484 20417
rect 20168 20451 20220 20460
rect 20168 20417 20177 20451
rect 20177 20417 20211 20451
rect 20211 20417 20220 20451
rect 20168 20408 20220 20417
rect 19524 20383 19576 20392
rect 19524 20349 19533 20383
rect 19533 20349 19567 20383
rect 19567 20349 19576 20383
rect 19524 20340 19576 20349
rect 19340 20272 19392 20324
rect 19708 20204 19760 20256
rect 20720 20451 20772 20460
rect 20720 20417 20729 20451
rect 20729 20417 20763 20451
rect 20763 20417 20772 20451
rect 20720 20408 20772 20417
rect 38292 20272 38344 20324
rect 37280 20204 37332 20256
rect 1950 20102 2002 20154
rect 2014 20102 2066 20154
rect 2078 20102 2130 20154
rect 2142 20102 2194 20154
rect 2206 20102 2258 20154
rect 6950 20102 7002 20154
rect 7014 20102 7066 20154
rect 7078 20102 7130 20154
rect 7142 20102 7194 20154
rect 7206 20102 7258 20154
rect 11950 20102 12002 20154
rect 12014 20102 12066 20154
rect 12078 20102 12130 20154
rect 12142 20102 12194 20154
rect 12206 20102 12258 20154
rect 16950 20102 17002 20154
rect 17014 20102 17066 20154
rect 17078 20102 17130 20154
rect 17142 20102 17194 20154
rect 17206 20102 17258 20154
rect 21950 20102 22002 20154
rect 22014 20102 22066 20154
rect 22078 20102 22130 20154
rect 22142 20102 22194 20154
rect 22206 20102 22258 20154
rect 26950 20102 27002 20154
rect 27014 20102 27066 20154
rect 27078 20102 27130 20154
rect 27142 20102 27194 20154
rect 27206 20102 27258 20154
rect 31950 20102 32002 20154
rect 32014 20102 32066 20154
rect 32078 20102 32130 20154
rect 32142 20102 32194 20154
rect 32206 20102 32258 20154
rect 36950 20102 37002 20154
rect 37014 20102 37066 20154
rect 37078 20102 37130 20154
rect 37142 20102 37194 20154
rect 37206 20102 37258 20154
rect 19524 19932 19576 19984
rect 19892 19932 19944 19984
rect 34520 19932 34572 19984
rect 38844 19932 38896 19984
rect 19800 19864 19852 19916
rect 940 19796 992 19848
rect 15292 19796 15344 19848
rect 22284 19796 22336 19848
rect 26240 19796 26292 19848
rect 19524 19728 19576 19780
rect 21732 19771 21784 19780
rect 21732 19737 21741 19771
rect 21741 19737 21775 19771
rect 21775 19737 21784 19771
rect 21732 19728 21784 19737
rect 18604 19703 18656 19712
rect 18604 19669 18613 19703
rect 18613 19669 18647 19703
rect 18647 19669 18656 19703
rect 18604 19660 18656 19669
rect 19708 19660 19760 19712
rect 20444 19703 20496 19712
rect 20444 19669 20453 19703
rect 20453 19669 20487 19703
rect 20487 19669 20496 19703
rect 20444 19660 20496 19669
rect 37280 19660 37332 19712
rect 2610 19558 2662 19610
rect 2674 19558 2726 19610
rect 2738 19558 2790 19610
rect 2802 19558 2854 19610
rect 2866 19558 2918 19610
rect 7610 19558 7662 19610
rect 7674 19558 7726 19610
rect 7738 19558 7790 19610
rect 7802 19558 7854 19610
rect 7866 19558 7918 19610
rect 12610 19558 12662 19610
rect 12674 19558 12726 19610
rect 12738 19558 12790 19610
rect 12802 19558 12854 19610
rect 12866 19558 12918 19610
rect 17610 19558 17662 19610
rect 17674 19558 17726 19610
rect 17738 19558 17790 19610
rect 17802 19558 17854 19610
rect 17866 19558 17918 19610
rect 22610 19558 22662 19610
rect 22674 19558 22726 19610
rect 22738 19558 22790 19610
rect 22802 19558 22854 19610
rect 22866 19558 22918 19610
rect 27610 19558 27662 19610
rect 27674 19558 27726 19610
rect 27738 19558 27790 19610
rect 27802 19558 27854 19610
rect 27866 19558 27918 19610
rect 32610 19558 32662 19610
rect 32674 19558 32726 19610
rect 32738 19558 32790 19610
rect 32802 19558 32854 19610
rect 32866 19558 32918 19610
rect 37610 19558 37662 19610
rect 37674 19558 37726 19610
rect 37738 19558 37790 19610
rect 37802 19558 37854 19610
rect 37866 19558 37918 19610
rect 18972 19499 19024 19508
rect 18972 19465 18981 19499
rect 18981 19465 19015 19499
rect 19015 19465 19024 19499
rect 18972 19456 19024 19465
rect 19340 19320 19392 19372
rect 21732 19456 21784 19508
rect 31760 19456 31812 19508
rect 26240 19388 26292 19440
rect 19708 19363 19760 19372
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 19892 19363 19944 19372
rect 19892 19329 19901 19363
rect 19901 19329 19935 19363
rect 19935 19329 19944 19363
rect 19892 19320 19944 19329
rect 20168 19363 20220 19372
rect 20168 19329 20177 19363
rect 20177 19329 20211 19363
rect 20211 19329 20220 19363
rect 20168 19320 20220 19329
rect 21088 19363 21140 19372
rect 21088 19329 21097 19363
rect 21097 19329 21131 19363
rect 21131 19329 21140 19363
rect 21088 19320 21140 19329
rect 38292 19363 38344 19372
rect 38292 19329 38301 19363
rect 38301 19329 38335 19363
rect 38335 19329 38344 19363
rect 38292 19320 38344 19329
rect 19800 19184 19852 19236
rect 1400 19159 1452 19168
rect 1400 19125 1409 19159
rect 1409 19125 1443 19159
rect 1443 19125 1452 19159
rect 1400 19116 1452 19125
rect 19524 19116 19576 19168
rect 20168 19116 20220 19168
rect 20352 19116 20404 19168
rect 20628 19184 20680 19236
rect 38476 19159 38528 19168
rect 38476 19125 38485 19159
rect 38485 19125 38519 19159
rect 38519 19125 38528 19159
rect 38476 19116 38528 19125
rect 1950 19014 2002 19066
rect 2014 19014 2066 19066
rect 2078 19014 2130 19066
rect 2142 19014 2194 19066
rect 2206 19014 2258 19066
rect 6950 19014 7002 19066
rect 7014 19014 7066 19066
rect 7078 19014 7130 19066
rect 7142 19014 7194 19066
rect 7206 19014 7258 19066
rect 11950 19014 12002 19066
rect 12014 19014 12066 19066
rect 12078 19014 12130 19066
rect 12142 19014 12194 19066
rect 12206 19014 12258 19066
rect 16950 19014 17002 19066
rect 17014 19014 17066 19066
rect 17078 19014 17130 19066
rect 17142 19014 17194 19066
rect 17206 19014 17258 19066
rect 21950 19014 22002 19066
rect 22014 19014 22066 19066
rect 22078 19014 22130 19066
rect 22142 19014 22194 19066
rect 22206 19014 22258 19066
rect 26950 19014 27002 19066
rect 27014 19014 27066 19066
rect 27078 19014 27130 19066
rect 27142 19014 27194 19066
rect 27206 19014 27258 19066
rect 31950 19014 32002 19066
rect 32014 19014 32066 19066
rect 32078 19014 32130 19066
rect 32142 19014 32194 19066
rect 32206 19014 32258 19066
rect 36950 19014 37002 19066
rect 37014 19014 37066 19066
rect 37078 19014 37130 19066
rect 37142 19014 37194 19066
rect 37206 19014 37258 19066
rect 22284 18912 22336 18964
rect 18604 18844 18656 18896
rect 19432 18776 19484 18828
rect 20444 18776 20496 18828
rect 940 18708 992 18760
rect 19524 18751 19576 18760
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 19708 18640 19760 18692
rect 19892 18572 19944 18624
rect 20352 18640 20404 18692
rect 20628 18615 20680 18624
rect 20628 18581 20637 18615
rect 20637 18581 20671 18615
rect 20671 18581 20680 18615
rect 20628 18572 20680 18581
rect 37280 18708 37332 18760
rect 21088 18572 21140 18624
rect 38476 18615 38528 18624
rect 38476 18581 38485 18615
rect 38485 18581 38519 18615
rect 38519 18581 38528 18615
rect 38476 18572 38528 18581
rect 2610 18470 2662 18522
rect 2674 18470 2726 18522
rect 2738 18470 2790 18522
rect 2802 18470 2854 18522
rect 2866 18470 2918 18522
rect 7610 18470 7662 18522
rect 7674 18470 7726 18522
rect 7738 18470 7790 18522
rect 7802 18470 7854 18522
rect 7866 18470 7918 18522
rect 12610 18470 12662 18522
rect 12674 18470 12726 18522
rect 12738 18470 12790 18522
rect 12802 18470 12854 18522
rect 12866 18470 12918 18522
rect 17610 18470 17662 18522
rect 17674 18470 17726 18522
rect 17738 18470 17790 18522
rect 17802 18470 17854 18522
rect 17866 18470 17918 18522
rect 22610 18470 22662 18522
rect 22674 18470 22726 18522
rect 22738 18470 22790 18522
rect 22802 18470 22854 18522
rect 22866 18470 22918 18522
rect 27610 18470 27662 18522
rect 27674 18470 27726 18522
rect 27738 18470 27790 18522
rect 27802 18470 27854 18522
rect 27866 18470 27918 18522
rect 32610 18470 32662 18522
rect 32674 18470 32726 18522
rect 32738 18470 32790 18522
rect 32802 18470 32854 18522
rect 32866 18470 32918 18522
rect 37610 18470 37662 18522
rect 37674 18470 37726 18522
rect 37738 18470 37790 18522
rect 37802 18470 37854 18522
rect 37866 18470 37918 18522
rect 19708 18368 19760 18420
rect 20720 18368 20772 18420
rect 19524 18343 19576 18352
rect 19524 18309 19533 18343
rect 19533 18309 19567 18343
rect 19567 18309 19576 18343
rect 19524 18300 19576 18309
rect 21088 18300 21140 18352
rect 19892 18232 19944 18284
rect 20628 18232 20680 18284
rect 1950 17926 2002 17978
rect 2014 17926 2066 17978
rect 2078 17926 2130 17978
rect 2142 17926 2194 17978
rect 2206 17926 2258 17978
rect 6950 17926 7002 17978
rect 7014 17926 7066 17978
rect 7078 17926 7130 17978
rect 7142 17926 7194 17978
rect 7206 17926 7258 17978
rect 11950 17926 12002 17978
rect 12014 17926 12066 17978
rect 12078 17926 12130 17978
rect 12142 17926 12194 17978
rect 12206 17926 12258 17978
rect 16950 17926 17002 17978
rect 17014 17926 17066 17978
rect 17078 17926 17130 17978
rect 17142 17926 17194 17978
rect 17206 17926 17258 17978
rect 21950 17926 22002 17978
rect 22014 17926 22066 17978
rect 22078 17926 22130 17978
rect 22142 17926 22194 17978
rect 22206 17926 22258 17978
rect 26950 17926 27002 17978
rect 27014 17926 27066 17978
rect 27078 17926 27130 17978
rect 27142 17926 27194 17978
rect 27206 17926 27258 17978
rect 31950 17926 32002 17978
rect 32014 17926 32066 17978
rect 32078 17926 32130 17978
rect 32142 17926 32194 17978
rect 32206 17926 32258 17978
rect 36950 17926 37002 17978
rect 37014 17926 37066 17978
rect 37078 17926 37130 17978
rect 37142 17926 37194 17978
rect 37206 17926 37258 17978
rect 31760 17824 31812 17876
rect 34520 17824 34572 17876
rect 2610 17382 2662 17434
rect 2674 17382 2726 17434
rect 2738 17382 2790 17434
rect 2802 17382 2854 17434
rect 2866 17382 2918 17434
rect 7610 17382 7662 17434
rect 7674 17382 7726 17434
rect 7738 17382 7790 17434
rect 7802 17382 7854 17434
rect 7866 17382 7918 17434
rect 12610 17382 12662 17434
rect 12674 17382 12726 17434
rect 12738 17382 12790 17434
rect 12802 17382 12854 17434
rect 12866 17382 12918 17434
rect 17610 17382 17662 17434
rect 17674 17382 17726 17434
rect 17738 17382 17790 17434
rect 17802 17382 17854 17434
rect 17866 17382 17918 17434
rect 22610 17382 22662 17434
rect 22674 17382 22726 17434
rect 22738 17382 22790 17434
rect 22802 17382 22854 17434
rect 22866 17382 22918 17434
rect 27610 17382 27662 17434
rect 27674 17382 27726 17434
rect 27738 17382 27790 17434
rect 27802 17382 27854 17434
rect 27866 17382 27918 17434
rect 32610 17382 32662 17434
rect 32674 17382 32726 17434
rect 32738 17382 32790 17434
rect 32802 17382 32854 17434
rect 32866 17382 32918 17434
rect 37610 17382 37662 17434
rect 37674 17382 37726 17434
rect 37738 17382 37790 17434
rect 37802 17382 37854 17434
rect 37866 17382 37918 17434
rect 1950 16838 2002 16890
rect 2014 16838 2066 16890
rect 2078 16838 2130 16890
rect 2142 16838 2194 16890
rect 2206 16838 2258 16890
rect 6950 16838 7002 16890
rect 7014 16838 7066 16890
rect 7078 16838 7130 16890
rect 7142 16838 7194 16890
rect 7206 16838 7258 16890
rect 11950 16838 12002 16890
rect 12014 16838 12066 16890
rect 12078 16838 12130 16890
rect 12142 16838 12194 16890
rect 12206 16838 12258 16890
rect 16950 16838 17002 16890
rect 17014 16838 17066 16890
rect 17078 16838 17130 16890
rect 17142 16838 17194 16890
rect 17206 16838 17258 16890
rect 21950 16838 22002 16890
rect 22014 16838 22066 16890
rect 22078 16838 22130 16890
rect 22142 16838 22194 16890
rect 22206 16838 22258 16890
rect 26950 16838 27002 16890
rect 27014 16838 27066 16890
rect 27078 16838 27130 16890
rect 27142 16838 27194 16890
rect 27206 16838 27258 16890
rect 31950 16838 32002 16890
rect 32014 16838 32066 16890
rect 32078 16838 32130 16890
rect 32142 16838 32194 16890
rect 32206 16838 32258 16890
rect 36950 16838 37002 16890
rect 37014 16838 37066 16890
rect 37078 16838 37130 16890
rect 37142 16838 37194 16890
rect 37206 16838 37258 16890
rect 2610 16294 2662 16346
rect 2674 16294 2726 16346
rect 2738 16294 2790 16346
rect 2802 16294 2854 16346
rect 2866 16294 2918 16346
rect 7610 16294 7662 16346
rect 7674 16294 7726 16346
rect 7738 16294 7790 16346
rect 7802 16294 7854 16346
rect 7866 16294 7918 16346
rect 12610 16294 12662 16346
rect 12674 16294 12726 16346
rect 12738 16294 12790 16346
rect 12802 16294 12854 16346
rect 12866 16294 12918 16346
rect 17610 16294 17662 16346
rect 17674 16294 17726 16346
rect 17738 16294 17790 16346
rect 17802 16294 17854 16346
rect 17866 16294 17918 16346
rect 22610 16294 22662 16346
rect 22674 16294 22726 16346
rect 22738 16294 22790 16346
rect 22802 16294 22854 16346
rect 22866 16294 22918 16346
rect 27610 16294 27662 16346
rect 27674 16294 27726 16346
rect 27738 16294 27790 16346
rect 27802 16294 27854 16346
rect 27866 16294 27918 16346
rect 32610 16294 32662 16346
rect 32674 16294 32726 16346
rect 32738 16294 32790 16346
rect 32802 16294 32854 16346
rect 32866 16294 32918 16346
rect 37610 16294 37662 16346
rect 37674 16294 37726 16346
rect 37738 16294 37790 16346
rect 37802 16294 37854 16346
rect 37866 16294 37918 16346
rect 1950 15750 2002 15802
rect 2014 15750 2066 15802
rect 2078 15750 2130 15802
rect 2142 15750 2194 15802
rect 2206 15750 2258 15802
rect 6950 15750 7002 15802
rect 7014 15750 7066 15802
rect 7078 15750 7130 15802
rect 7142 15750 7194 15802
rect 7206 15750 7258 15802
rect 11950 15750 12002 15802
rect 12014 15750 12066 15802
rect 12078 15750 12130 15802
rect 12142 15750 12194 15802
rect 12206 15750 12258 15802
rect 16950 15750 17002 15802
rect 17014 15750 17066 15802
rect 17078 15750 17130 15802
rect 17142 15750 17194 15802
rect 17206 15750 17258 15802
rect 21950 15750 22002 15802
rect 22014 15750 22066 15802
rect 22078 15750 22130 15802
rect 22142 15750 22194 15802
rect 22206 15750 22258 15802
rect 26950 15750 27002 15802
rect 27014 15750 27066 15802
rect 27078 15750 27130 15802
rect 27142 15750 27194 15802
rect 27206 15750 27258 15802
rect 31950 15750 32002 15802
rect 32014 15750 32066 15802
rect 32078 15750 32130 15802
rect 32142 15750 32194 15802
rect 32206 15750 32258 15802
rect 36950 15750 37002 15802
rect 37014 15750 37066 15802
rect 37078 15750 37130 15802
rect 37142 15750 37194 15802
rect 37206 15750 37258 15802
rect 2610 15206 2662 15258
rect 2674 15206 2726 15258
rect 2738 15206 2790 15258
rect 2802 15206 2854 15258
rect 2866 15206 2918 15258
rect 7610 15206 7662 15258
rect 7674 15206 7726 15258
rect 7738 15206 7790 15258
rect 7802 15206 7854 15258
rect 7866 15206 7918 15258
rect 12610 15206 12662 15258
rect 12674 15206 12726 15258
rect 12738 15206 12790 15258
rect 12802 15206 12854 15258
rect 12866 15206 12918 15258
rect 17610 15206 17662 15258
rect 17674 15206 17726 15258
rect 17738 15206 17790 15258
rect 17802 15206 17854 15258
rect 17866 15206 17918 15258
rect 22610 15206 22662 15258
rect 22674 15206 22726 15258
rect 22738 15206 22790 15258
rect 22802 15206 22854 15258
rect 22866 15206 22918 15258
rect 27610 15206 27662 15258
rect 27674 15206 27726 15258
rect 27738 15206 27790 15258
rect 27802 15206 27854 15258
rect 27866 15206 27918 15258
rect 32610 15206 32662 15258
rect 32674 15206 32726 15258
rect 32738 15206 32790 15258
rect 32802 15206 32854 15258
rect 32866 15206 32918 15258
rect 37610 15206 37662 15258
rect 37674 15206 37726 15258
rect 37738 15206 37790 15258
rect 37802 15206 37854 15258
rect 37866 15206 37918 15258
rect 1950 14662 2002 14714
rect 2014 14662 2066 14714
rect 2078 14662 2130 14714
rect 2142 14662 2194 14714
rect 2206 14662 2258 14714
rect 6950 14662 7002 14714
rect 7014 14662 7066 14714
rect 7078 14662 7130 14714
rect 7142 14662 7194 14714
rect 7206 14662 7258 14714
rect 11950 14662 12002 14714
rect 12014 14662 12066 14714
rect 12078 14662 12130 14714
rect 12142 14662 12194 14714
rect 12206 14662 12258 14714
rect 16950 14662 17002 14714
rect 17014 14662 17066 14714
rect 17078 14662 17130 14714
rect 17142 14662 17194 14714
rect 17206 14662 17258 14714
rect 21950 14662 22002 14714
rect 22014 14662 22066 14714
rect 22078 14662 22130 14714
rect 22142 14662 22194 14714
rect 22206 14662 22258 14714
rect 26950 14662 27002 14714
rect 27014 14662 27066 14714
rect 27078 14662 27130 14714
rect 27142 14662 27194 14714
rect 27206 14662 27258 14714
rect 31950 14662 32002 14714
rect 32014 14662 32066 14714
rect 32078 14662 32130 14714
rect 32142 14662 32194 14714
rect 32206 14662 32258 14714
rect 36950 14662 37002 14714
rect 37014 14662 37066 14714
rect 37078 14662 37130 14714
rect 37142 14662 37194 14714
rect 37206 14662 37258 14714
rect 2610 14118 2662 14170
rect 2674 14118 2726 14170
rect 2738 14118 2790 14170
rect 2802 14118 2854 14170
rect 2866 14118 2918 14170
rect 7610 14118 7662 14170
rect 7674 14118 7726 14170
rect 7738 14118 7790 14170
rect 7802 14118 7854 14170
rect 7866 14118 7918 14170
rect 12610 14118 12662 14170
rect 12674 14118 12726 14170
rect 12738 14118 12790 14170
rect 12802 14118 12854 14170
rect 12866 14118 12918 14170
rect 17610 14118 17662 14170
rect 17674 14118 17726 14170
rect 17738 14118 17790 14170
rect 17802 14118 17854 14170
rect 17866 14118 17918 14170
rect 22610 14118 22662 14170
rect 22674 14118 22726 14170
rect 22738 14118 22790 14170
rect 22802 14118 22854 14170
rect 22866 14118 22918 14170
rect 27610 14118 27662 14170
rect 27674 14118 27726 14170
rect 27738 14118 27790 14170
rect 27802 14118 27854 14170
rect 27866 14118 27918 14170
rect 32610 14118 32662 14170
rect 32674 14118 32726 14170
rect 32738 14118 32790 14170
rect 32802 14118 32854 14170
rect 32866 14118 32918 14170
rect 37610 14118 37662 14170
rect 37674 14118 37726 14170
rect 37738 14118 37790 14170
rect 37802 14118 37854 14170
rect 37866 14118 37918 14170
rect 1950 13574 2002 13626
rect 2014 13574 2066 13626
rect 2078 13574 2130 13626
rect 2142 13574 2194 13626
rect 2206 13574 2258 13626
rect 6950 13574 7002 13626
rect 7014 13574 7066 13626
rect 7078 13574 7130 13626
rect 7142 13574 7194 13626
rect 7206 13574 7258 13626
rect 11950 13574 12002 13626
rect 12014 13574 12066 13626
rect 12078 13574 12130 13626
rect 12142 13574 12194 13626
rect 12206 13574 12258 13626
rect 16950 13574 17002 13626
rect 17014 13574 17066 13626
rect 17078 13574 17130 13626
rect 17142 13574 17194 13626
rect 17206 13574 17258 13626
rect 21950 13574 22002 13626
rect 22014 13574 22066 13626
rect 22078 13574 22130 13626
rect 22142 13574 22194 13626
rect 22206 13574 22258 13626
rect 26950 13574 27002 13626
rect 27014 13574 27066 13626
rect 27078 13574 27130 13626
rect 27142 13574 27194 13626
rect 27206 13574 27258 13626
rect 31950 13574 32002 13626
rect 32014 13574 32066 13626
rect 32078 13574 32130 13626
rect 32142 13574 32194 13626
rect 32206 13574 32258 13626
rect 36950 13574 37002 13626
rect 37014 13574 37066 13626
rect 37078 13574 37130 13626
rect 37142 13574 37194 13626
rect 37206 13574 37258 13626
rect 2610 13030 2662 13082
rect 2674 13030 2726 13082
rect 2738 13030 2790 13082
rect 2802 13030 2854 13082
rect 2866 13030 2918 13082
rect 7610 13030 7662 13082
rect 7674 13030 7726 13082
rect 7738 13030 7790 13082
rect 7802 13030 7854 13082
rect 7866 13030 7918 13082
rect 12610 13030 12662 13082
rect 12674 13030 12726 13082
rect 12738 13030 12790 13082
rect 12802 13030 12854 13082
rect 12866 13030 12918 13082
rect 17610 13030 17662 13082
rect 17674 13030 17726 13082
rect 17738 13030 17790 13082
rect 17802 13030 17854 13082
rect 17866 13030 17918 13082
rect 22610 13030 22662 13082
rect 22674 13030 22726 13082
rect 22738 13030 22790 13082
rect 22802 13030 22854 13082
rect 22866 13030 22918 13082
rect 27610 13030 27662 13082
rect 27674 13030 27726 13082
rect 27738 13030 27790 13082
rect 27802 13030 27854 13082
rect 27866 13030 27918 13082
rect 32610 13030 32662 13082
rect 32674 13030 32726 13082
rect 32738 13030 32790 13082
rect 32802 13030 32854 13082
rect 32866 13030 32918 13082
rect 37610 13030 37662 13082
rect 37674 13030 37726 13082
rect 37738 13030 37790 13082
rect 37802 13030 37854 13082
rect 37866 13030 37918 13082
rect 1950 12486 2002 12538
rect 2014 12486 2066 12538
rect 2078 12486 2130 12538
rect 2142 12486 2194 12538
rect 2206 12486 2258 12538
rect 6950 12486 7002 12538
rect 7014 12486 7066 12538
rect 7078 12486 7130 12538
rect 7142 12486 7194 12538
rect 7206 12486 7258 12538
rect 11950 12486 12002 12538
rect 12014 12486 12066 12538
rect 12078 12486 12130 12538
rect 12142 12486 12194 12538
rect 12206 12486 12258 12538
rect 16950 12486 17002 12538
rect 17014 12486 17066 12538
rect 17078 12486 17130 12538
rect 17142 12486 17194 12538
rect 17206 12486 17258 12538
rect 21950 12486 22002 12538
rect 22014 12486 22066 12538
rect 22078 12486 22130 12538
rect 22142 12486 22194 12538
rect 22206 12486 22258 12538
rect 26950 12486 27002 12538
rect 27014 12486 27066 12538
rect 27078 12486 27130 12538
rect 27142 12486 27194 12538
rect 27206 12486 27258 12538
rect 31950 12486 32002 12538
rect 32014 12486 32066 12538
rect 32078 12486 32130 12538
rect 32142 12486 32194 12538
rect 32206 12486 32258 12538
rect 36950 12486 37002 12538
rect 37014 12486 37066 12538
rect 37078 12486 37130 12538
rect 37142 12486 37194 12538
rect 37206 12486 37258 12538
rect 2610 11942 2662 11994
rect 2674 11942 2726 11994
rect 2738 11942 2790 11994
rect 2802 11942 2854 11994
rect 2866 11942 2918 11994
rect 7610 11942 7662 11994
rect 7674 11942 7726 11994
rect 7738 11942 7790 11994
rect 7802 11942 7854 11994
rect 7866 11942 7918 11994
rect 12610 11942 12662 11994
rect 12674 11942 12726 11994
rect 12738 11942 12790 11994
rect 12802 11942 12854 11994
rect 12866 11942 12918 11994
rect 17610 11942 17662 11994
rect 17674 11942 17726 11994
rect 17738 11942 17790 11994
rect 17802 11942 17854 11994
rect 17866 11942 17918 11994
rect 22610 11942 22662 11994
rect 22674 11942 22726 11994
rect 22738 11942 22790 11994
rect 22802 11942 22854 11994
rect 22866 11942 22918 11994
rect 27610 11942 27662 11994
rect 27674 11942 27726 11994
rect 27738 11942 27790 11994
rect 27802 11942 27854 11994
rect 27866 11942 27918 11994
rect 32610 11942 32662 11994
rect 32674 11942 32726 11994
rect 32738 11942 32790 11994
rect 32802 11942 32854 11994
rect 32866 11942 32918 11994
rect 37610 11942 37662 11994
rect 37674 11942 37726 11994
rect 37738 11942 37790 11994
rect 37802 11942 37854 11994
rect 37866 11942 37918 11994
rect 1950 11398 2002 11450
rect 2014 11398 2066 11450
rect 2078 11398 2130 11450
rect 2142 11398 2194 11450
rect 2206 11398 2258 11450
rect 6950 11398 7002 11450
rect 7014 11398 7066 11450
rect 7078 11398 7130 11450
rect 7142 11398 7194 11450
rect 7206 11398 7258 11450
rect 11950 11398 12002 11450
rect 12014 11398 12066 11450
rect 12078 11398 12130 11450
rect 12142 11398 12194 11450
rect 12206 11398 12258 11450
rect 16950 11398 17002 11450
rect 17014 11398 17066 11450
rect 17078 11398 17130 11450
rect 17142 11398 17194 11450
rect 17206 11398 17258 11450
rect 21950 11398 22002 11450
rect 22014 11398 22066 11450
rect 22078 11398 22130 11450
rect 22142 11398 22194 11450
rect 22206 11398 22258 11450
rect 26950 11398 27002 11450
rect 27014 11398 27066 11450
rect 27078 11398 27130 11450
rect 27142 11398 27194 11450
rect 27206 11398 27258 11450
rect 31950 11398 32002 11450
rect 32014 11398 32066 11450
rect 32078 11398 32130 11450
rect 32142 11398 32194 11450
rect 32206 11398 32258 11450
rect 36950 11398 37002 11450
rect 37014 11398 37066 11450
rect 37078 11398 37130 11450
rect 37142 11398 37194 11450
rect 37206 11398 37258 11450
rect 2610 10854 2662 10906
rect 2674 10854 2726 10906
rect 2738 10854 2790 10906
rect 2802 10854 2854 10906
rect 2866 10854 2918 10906
rect 7610 10854 7662 10906
rect 7674 10854 7726 10906
rect 7738 10854 7790 10906
rect 7802 10854 7854 10906
rect 7866 10854 7918 10906
rect 12610 10854 12662 10906
rect 12674 10854 12726 10906
rect 12738 10854 12790 10906
rect 12802 10854 12854 10906
rect 12866 10854 12918 10906
rect 17610 10854 17662 10906
rect 17674 10854 17726 10906
rect 17738 10854 17790 10906
rect 17802 10854 17854 10906
rect 17866 10854 17918 10906
rect 22610 10854 22662 10906
rect 22674 10854 22726 10906
rect 22738 10854 22790 10906
rect 22802 10854 22854 10906
rect 22866 10854 22918 10906
rect 27610 10854 27662 10906
rect 27674 10854 27726 10906
rect 27738 10854 27790 10906
rect 27802 10854 27854 10906
rect 27866 10854 27918 10906
rect 32610 10854 32662 10906
rect 32674 10854 32726 10906
rect 32738 10854 32790 10906
rect 32802 10854 32854 10906
rect 32866 10854 32918 10906
rect 37610 10854 37662 10906
rect 37674 10854 37726 10906
rect 37738 10854 37790 10906
rect 37802 10854 37854 10906
rect 37866 10854 37918 10906
rect 1950 10310 2002 10362
rect 2014 10310 2066 10362
rect 2078 10310 2130 10362
rect 2142 10310 2194 10362
rect 2206 10310 2258 10362
rect 6950 10310 7002 10362
rect 7014 10310 7066 10362
rect 7078 10310 7130 10362
rect 7142 10310 7194 10362
rect 7206 10310 7258 10362
rect 11950 10310 12002 10362
rect 12014 10310 12066 10362
rect 12078 10310 12130 10362
rect 12142 10310 12194 10362
rect 12206 10310 12258 10362
rect 16950 10310 17002 10362
rect 17014 10310 17066 10362
rect 17078 10310 17130 10362
rect 17142 10310 17194 10362
rect 17206 10310 17258 10362
rect 21950 10310 22002 10362
rect 22014 10310 22066 10362
rect 22078 10310 22130 10362
rect 22142 10310 22194 10362
rect 22206 10310 22258 10362
rect 26950 10310 27002 10362
rect 27014 10310 27066 10362
rect 27078 10310 27130 10362
rect 27142 10310 27194 10362
rect 27206 10310 27258 10362
rect 31950 10310 32002 10362
rect 32014 10310 32066 10362
rect 32078 10310 32130 10362
rect 32142 10310 32194 10362
rect 32206 10310 32258 10362
rect 36950 10310 37002 10362
rect 37014 10310 37066 10362
rect 37078 10310 37130 10362
rect 37142 10310 37194 10362
rect 37206 10310 37258 10362
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 7610 9766 7662 9818
rect 7674 9766 7726 9818
rect 7738 9766 7790 9818
rect 7802 9766 7854 9818
rect 7866 9766 7918 9818
rect 12610 9766 12662 9818
rect 12674 9766 12726 9818
rect 12738 9766 12790 9818
rect 12802 9766 12854 9818
rect 12866 9766 12918 9818
rect 17610 9766 17662 9818
rect 17674 9766 17726 9818
rect 17738 9766 17790 9818
rect 17802 9766 17854 9818
rect 17866 9766 17918 9818
rect 22610 9766 22662 9818
rect 22674 9766 22726 9818
rect 22738 9766 22790 9818
rect 22802 9766 22854 9818
rect 22866 9766 22918 9818
rect 27610 9766 27662 9818
rect 27674 9766 27726 9818
rect 27738 9766 27790 9818
rect 27802 9766 27854 9818
rect 27866 9766 27918 9818
rect 32610 9766 32662 9818
rect 32674 9766 32726 9818
rect 32738 9766 32790 9818
rect 32802 9766 32854 9818
rect 32866 9766 32918 9818
rect 37610 9766 37662 9818
rect 37674 9766 37726 9818
rect 37738 9766 37790 9818
rect 37802 9766 37854 9818
rect 37866 9766 37918 9818
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6950 9222 7002 9274
rect 7014 9222 7066 9274
rect 7078 9222 7130 9274
rect 7142 9222 7194 9274
rect 7206 9222 7258 9274
rect 11950 9222 12002 9274
rect 12014 9222 12066 9274
rect 12078 9222 12130 9274
rect 12142 9222 12194 9274
rect 12206 9222 12258 9274
rect 16950 9222 17002 9274
rect 17014 9222 17066 9274
rect 17078 9222 17130 9274
rect 17142 9222 17194 9274
rect 17206 9222 17258 9274
rect 21950 9222 22002 9274
rect 22014 9222 22066 9274
rect 22078 9222 22130 9274
rect 22142 9222 22194 9274
rect 22206 9222 22258 9274
rect 26950 9222 27002 9274
rect 27014 9222 27066 9274
rect 27078 9222 27130 9274
rect 27142 9222 27194 9274
rect 27206 9222 27258 9274
rect 31950 9222 32002 9274
rect 32014 9222 32066 9274
rect 32078 9222 32130 9274
rect 32142 9222 32194 9274
rect 32206 9222 32258 9274
rect 36950 9222 37002 9274
rect 37014 9222 37066 9274
rect 37078 9222 37130 9274
rect 37142 9222 37194 9274
rect 37206 9222 37258 9274
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 7610 8678 7662 8730
rect 7674 8678 7726 8730
rect 7738 8678 7790 8730
rect 7802 8678 7854 8730
rect 7866 8678 7918 8730
rect 12610 8678 12662 8730
rect 12674 8678 12726 8730
rect 12738 8678 12790 8730
rect 12802 8678 12854 8730
rect 12866 8678 12918 8730
rect 17610 8678 17662 8730
rect 17674 8678 17726 8730
rect 17738 8678 17790 8730
rect 17802 8678 17854 8730
rect 17866 8678 17918 8730
rect 22610 8678 22662 8730
rect 22674 8678 22726 8730
rect 22738 8678 22790 8730
rect 22802 8678 22854 8730
rect 22866 8678 22918 8730
rect 27610 8678 27662 8730
rect 27674 8678 27726 8730
rect 27738 8678 27790 8730
rect 27802 8678 27854 8730
rect 27866 8678 27918 8730
rect 32610 8678 32662 8730
rect 32674 8678 32726 8730
rect 32738 8678 32790 8730
rect 32802 8678 32854 8730
rect 32866 8678 32918 8730
rect 37610 8678 37662 8730
rect 37674 8678 37726 8730
rect 37738 8678 37790 8730
rect 37802 8678 37854 8730
rect 37866 8678 37918 8730
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 6950 8134 7002 8186
rect 7014 8134 7066 8186
rect 7078 8134 7130 8186
rect 7142 8134 7194 8186
rect 7206 8134 7258 8186
rect 11950 8134 12002 8186
rect 12014 8134 12066 8186
rect 12078 8134 12130 8186
rect 12142 8134 12194 8186
rect 12206 8134 12258 8186
rect 16950 8134 17002 8186
rect 17014 8134 17066 8186
rect 17078 8134 17130 8186
rect 17142 8134 17194 8186
rect 17206 8134 17258 8186
rect 21950 8134 22002 8186
rect 22014 8134 22066 8186
rect 22078 8134 22130 8186
rect 22142 8134 22194 8186
rect 22206 8134 22258 8186
rect 26950 8134 27002 8186
rect 27014 8134 27066 8186
rect 27078 8134 27130 8186
rect 27142 8134 27194 8186
rect 27206 8134 27258 8186
rect 31950 8134 32002 8186
rect 32014 8134 32066 8186
rect 32078 8134 32130 8186
rect 32142 8134 32194 8186
rect 32206 8134 32258 8186
rect 36950 8134 37002 8186
rect 37014 8134 37066 8186
rect 37078 8134 37130 8186
rect 37142 8134 37194 8186
rect 37206 8134 37258 8186
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 7610 7590 7662 7642
rect 7674 7590 7726 7642
rect 7738 7590 7790 7642
rect 7802 7590 7854 7642
rect 7866 7590 7918 7642
rect 12610 7590 12662 7642
rect 12674 7590 12726 7642
rect 12738 7590 12790 7642
rect 12802 7590 12854 7642
rect 12866 7590 12918 7642
rect 17610 7590 17662 7642
rect 17674 7590 17726 7642
rect 17738 7590 17790 7642
rect 17802 7590 17854 7642
rect 17866 7590 17918 7642
rect 22610 7590 22662 7642
rect 22674 7590 22726 7642
rect 22738 7590 22790 7642
rect 22802 7590 22854 7642
rect 22866 7590 22918 7642
rect 27610 7590 27662 7642
rect 27674 7590 27726 7642
rect 27738 7590 27790 7642
rect 27802 7590 27854 7642
rect 27866 7590 27918 7642
rect 32610 7590 32662 7642
rect 32674 7590 32726 7642
rect 32738 7590 32790 7642
rect 32802 7590 32854 7642
rect 32866 7590 32918 7642
rect 37610 7590 37662 7642
rect 37674 7590 37726 7642
rect 37738 7590 37790 7642
rect 37802 7590 37854 7642
rect 37866 7590 37918 7642
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 6950 7046 7002 7098
rect 7014 7046 7066 7098
rect 7078 7046 7130 7098
rect 7142 7046 7194 7098
rect 7206 7046 7258 7098
rect 11950 7046 12002 7098
rect 12014 7046 12066 7098
rect 12078 7046 12130 7098
rect 12142 7046 12194 7098
rect 12206 7046 12258 7098
rect 16950 7046 17002 7098
rect 17014 7046 17066 7098
rect 17078 7046 17130 7098
rect 17142 7046 17194 7098
rect 17206 7046 17258 7098
rect 21950 7046 22002 7098
rect 22014 7046 22066 7098
rect 22078 7046 22130 7098
rect 22142 7046 22194 7098
rect 22206 7046 22258 7098
rect 26950 7046 27002 7098
rect 27014 7046 27066 7098
rect 27078 7046 27130 7098
rect 27142 7046 27194 7098
rect 27206 7046 27258 7098
rect 31950 7046 32002 7098
rect 32014 7046 32066 7098
rect 32078 7046 32130 7098
rect 32142 7046 32194 7098
rect 32206 7046 32258 7098
rect 36950 7046 37002 7098
rect 37014 7046 37066 7098
rect 37078 7046 37130 7098
rect 37142 7046 37194 7098
rect 37206 7046 37258 7098
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 7610 6502 7662 6554
rect 7674 6502 7726 6554
rect 7738 6502 7790 6554
rect 7802 6502 7854 6554
rect 7866 6502 7918 6554
rect 12610 6502 12662 6554
rect 12674 6502 12726 6554
rect 12738 6502 12790 6554
rect 12802 6502 12854 6554
rect 12866 6502 12918 6554
rect 17610 6502 17662 6554
rect 17674 6502 17726 6554
rect 17738 6502 17790 6554
rect 17802 6502 17854 6554
rect 17866 6502 17918 6554
rect 22610 6502 22662 6554
rect 22674 6502 22726 6554
rect 22738 6502 22790 6554
rect 22802 6502 22854 6554
rect 22866 6502 22918 6554
rect 27610 6502 27662 6554
rect 27674 6502 27726 6554
rect 27738 6502 27790 6554
rect 27802 6502 27854 6554
rect 27866 6502 27918 6554
rect 32610 6502 32662 6554
rect 32674 6502 32726 6554
rect 32738 6502 32790 6554
rect 32802 6502 32854 6554
rect 32866 6502 32918 6554
rect 37610 6502 37662 6554
rect 37674 6502 37726 6554
rect 37738 6502 37790 6554
rect 37802 6502 37854 6554
rect 37866 6502 37918 6554
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 6950 5958 7002 6010
rect 7014 5958 7066 6010
rect 7078 5958 7130 6010
rect 7142 5958 7194 6010
rect 7206 5958 7258 6010
rect 11950 5958 12002 6010
rect 12014 5958 12066 6010
rect 12078 5958 12130 6010
rect 12142 5958 12194 6010
rect 12206 5958 12258 6010
rect 16950 5958 17002 6010
rect 17014 5958 17066 6010
rect 17078 5958 17130 6010
rect 17142 5958 17194 6010
rect 17206 5958 17258 6010
rect 21950 5958 22002 6010
rect 22014 5958 22066 6010
rect 22078 5958 22130 6010
rect 22142 5958 22194 6010
rect 22206 5958 22258 6010
rect 26950 5958 27002 6010
rect 27014 5958 27066 6010
rect 27078 5958 27130 6010
rect 27142 5958 27194 6010
rect 27206 5958 27258 6010
rect 31950 5958 32002 6010
rect 32014 5958 32066 6010
rect 32078 5958 32130 6010
rect 32142 5958 32194 6010
rect 32206 5958 32258 6010
rect 36950 5958 37002 6010
rect 37014 5958 37066 6010
rect 37078 5958 37130 6010
rect 37142 5958 37194 6010
rect 37206 5958 37258 6010
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 7610 5414 7662 5466
rect 7674 5414 7726 5466
rect 7738 5414 7790 5466
rect 7802 5414 7854 5466
rect 7866 5414 7918 5466
rect 12610 5414 12662 5466
rect 12674 5414 12726 5466
rect 12738 5414 12790 5466
rect 12802 5414 12854 5466
rect 12866 5414 12918 5466
rect 17610 5414 17662 5466
rect 17674 5414 17726 5466
rect 17738 5414 17790 5466
rect 17802 5414 17854 5466
rect 17866 5414 17918 5466
rect 22610 5414 22662 5466
rect 22674 5414 22726 5466
rect 22738 5414 22790 5466
rect 22802 5414 22854 5466
rect 22866 5414 22918 5466
rect 27610 5414 27662 5466
rect 27674 5414 27726 5466
rect 27738 5414 27790 5466
rect 27802 5414 27854 5466
rect 27866 5414 27918 5466
rect 32610 5414 32662 5466
rect 32674 5414 32726 5466
rect 32738 5414 32790 5466
rect 32802 5414 32854 5466
rect 32866 5414 32918 5466
rect 37610 5414 37662 5466
rect 37674 5414 37726 5466
rect 37738 5414 37790 5466
rect 37802 5414 37854 5466
rect 37866 5414 37918 5466
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 6950 4870 7002 4922
rect 7014 4870 7066 4922
rect 7078 4870 7130 4922
rect 7142 4870 7194 4922
rect 7206 4870 7258 4922
rect 11950 4870 12002 4922
rect 12014 4870 12066 4922
rect 12078 4870 12130 4922
rect 12142 4870 12194 4922
rect 12206 4870 12258 4922
rect 16950 4870 17002 4922
rect 17014 4870 17066 4922
rect 17078 4870 17130 4922
rect 17142 4870 17194 4922
rect 17206 4870 17258 4922
rect 21950 4870 22002 4922
rect 22014 4870 22066 4922
rect 22078 4870 22130 4922
rect 22142 4870 22194 4922
rect 22206 4870 22258 4922
rect 26950 4870 27002 4922
rect 27014 4870 27066 4922
rect 27078 4870 27130 4922
rect 27142 4870 27194 4922
rect 27206 4870 27258 4922
rect 31950 4870 32002 4922
rect 32014 4870 32066 4922
rect 32078 4870 32130 4922
rect 32142 4870 32194 4922
rect 32206 4870 32258 4922
rect 36950 4870 37002 4922
rect 37014 4870 37066 4922
rect 37078 4870 37130 4922
rect 37142 4870 37194 4922
rect 37206 4870 37258 4922
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 7610 4326 7662 4378
rect 7674 4326 7726 4378
rect 7738 4326 7790 4378
rect 7802 4326 7854 4378
rect 7866 4326 7918 4378
rect 12610 4326 12662 4378
rect 12674 4326 12726 4378
rect 12738 4326 12790 4378
rect 12802 4326 12854 4378
rect 12866 4326 12918 4378
rect 17610 4326 17662 4378
rect 17674 4326 17726 4378
rect 17738 4326 17790 4378
rect 17802 4326 17854 4378
rect 17866 4326 17918 4378
rect 22610 4326 22662 4378
rect 22674 4326 22726 4378
rect 22738 4326 22790 4378
rect 22802 4326 22854 4378
rect 22866 4326 22918 4378
rect 27610 4326 27662 4378
rect 27674 4326 27726 4378
rect 27738 4326 27790 4378
rect 27802 4326 27854 4378
rect 27866 4326 27918 4378
rect 32610 4326 32662 4378
rect 32674 4326 32726 4378
rect 32738 4326 32790 4378
rect 32802 4326 32854 4378
rect 32866 4326 32918 4378
rect 37610 4326 37662 4378
rect 37674 4326 37726 4378
rect 37738 4326 37790 4378
rect 37802 4326 37854 4378
rect 37866 4326 37918 4378
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 6950 3782 7002 3834
rect 7014 3782 7066 3834
rect 7078 3782 7130 3834
rect 7142 3782 7194 3834
rect 7206 3782 7258 3834
rect 11950 3782 12002 3834
rect 12014 3782 12066 3834
rect 12078 3782 12130 3834
rect 12142 3782 12194 3834
rect 12206 3782 12258 3834
rect 16950 3782 17002 3834
rect 17014 3782 17066 3834
rect 17078 3782 17130 3834
rect 17142 3782 17194 3834
rect 17206 3782 17258 3834
rect 21950 3782 22002 3834
rect 22014 3782 22066 3834
rect 22078 3782 22130 3834
rect 22142 3782 22194 3834
rect 22206 3782 22258 3834
rect 26950 3782 27002 3834
rect 27014 3782 27066 3834
rect 27078 3782 27130 3834
rect 27142 3782 27194 3834
rect 27206 3782 27258 3834
rect 31950 3782 32002 3834
rect 32014 3782 32066 3834
rect 32078 3782 32130 3834
rect 32142 3782 32194 3834
rect 32206 3782 32258 3834
rect 36950 3782 37002 3834
rect 37014 3782 37066 3834
rect 37078 3782 37130 3834
rect 37142 3782 37194 3834
rect 37206 3782 37258 3834
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 7610 3238 7662 3290
rect 7674 3238 7726 3290
rect 7738 3238 7790 3290
rect 7802 3238 7854 3290
rect 7866 3238 7918 3290
rect 12610 3238 12662 3290
rect 12674 3238 12726 3290
rect 12738 3238 12790 3290
rect 12802 3238 12854 3290
rect 12866 3238 12918 3290
rect 17610 3238 17662 3290
rect 17674 3238 17726 3290
rect 17738 3238 17790 3290
rect 17802 3238 17854 3290
rect 17866 3238 17918 3290
rect 22610 3238 22662 3290
rect 22674 3238 22726 3290
rect 22738 3238 22790 3290
rect 22802 3238 22854 3290
rect 22866 3238 22918 3290
rect 27610 3238 27662 3290
rect 27674 3238 27726 3290
rect 27738 3238 27790 3290
rect 27802 3238 27854 3290
rect 27866 3238 27918 3290
rect 32610 3238 32662 3290
rect 32674 3238 32726 3290
rect 32738 3238 32790 3290
rect 32802 3238 32854 3290
rect 32866 3238 32918 3290
rect 37610 3238 37662 3290
rect 37674 3238 37726 3290
rect 37738 3238 37790 3290
rect 37802 3238 37854 3290
rect 37866 3238 37918 3290
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 6950 2694 7002 2746
rect 7014 2694 7066 2746
rect 7078 2694 7130 2746
rect 7142 2694 7194 2746
rect 7206 2694 7258 2746
rect 11950 2694 12002 2746
rect 12014 2694 12066 2746
rect 12078 2694 12130 2746
rect 12142 2694 12194 2746
rect 12206 2694 12258 2746
rect 16950 2694 17002 2746
rect 17014 2694 17066 2746
rect 17078 2694 17130 2746
rect 17142 2694 17194 2746
rect 17206 2694 17258 2746
rect 21950 2694 22002 2746
rect 22014 2694 22066 2746
rect 22078 2694 22130 2746
rect 22142 2694 22194 2746
rect 22206 2694 22258 2746
rect 26950 2694 27002 2746
rect 27014 2694 27066 2746
rect 27078 2694 27130 2746
rect 27142 2694 27194 2746
rect 27206 2694 27258 2746
rect 31950 2694 32002 2746
rect 32014 2694 32066 2746
rect 32078 2694 32130 2746
rect 32142 2694 32194 2746
rect 32206 2694 32258 2746
rect 36950 2694 37002 2746
rect 37014 2694 37066 2746
rect 37078 2694 37130 2746
rect 37142 2694 37194 2746
rect 37206 2694 37258 2746
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 7610 2150 7662 2202
rect 7674 2150 7726 2202
rect 7738 2150 7790 2202
rect 7802 2150 7854 2202
rect 7866 2150 7918 2202
rect 12610 2150 12662 2202
rect 12674 2150 12726 2202
rect 12738 2150 12790 2202
rect 12802 2150 12854 2202
rect 12866 2150 12918 2202
rect 17610 2150 17662 2202
rect 17674 2150 17726 2202
rect 17738 2150 17790 2202
rect 17802 2150 17854 2202
rect 17866 2150 17918 2202
rect 22610 2150 22662 2202
rect 22674 2150 22726 2202
rect 22738 2150 22790 2202
rect 22802 2150 22854 2202
rect 22866 2150 22918 2202
rect 27610 2150 27662 2202
rect 27674 2150 27726 2202
rect 27738 2150 27790 2202
rect 27802 2150 27854 2202
rect 27866 2150 27918 2202
rect 32610 2150 32662 2202
rect 32674 2150 32726 2202
rect 32738 2150 32790 2202
rect 32802 2150 32854 2202
rect 32866 2150 32918 2202
rect 37610 2150 37662 2202
rect 37674 2150 37726 2202
rect 37738 2150 37790 2202
rect 37802 2150 37854 2202
rect 37866 2150 37918 2202
<< metal2 >>
rect 1950 37564 2258 37573
rect 1950 37562 1956 37564
rect 2012 37562 2036 37564
rect 2092 37562 2116 37564
rect 2172 37562 2196 37564
rect 2252 37562 2258 37564
rect 2012 37510 2014 37562
rect 2194 37510 2196 37562
rect 1950 37508 1956 37510
rect 2012 37508 2036 37510
rect 2092 37508 2116 37510
rect 2172 37508 2196 37510
rect 2252 37508 2258 37510
rect 1950 37499 2258 37508
rect 6950 37564 7258 37573
rect 6950 37562 6956 37564
rect 7012 37562 7036 37564
rect 7092 37562 7116 37564
rect 7172 37562 7196 37564
rect 7252 37562 7258 37564
rect 7012 37510 7014 37562
rect 7194 37510 7196 37562
rect 6950 37508 6956 37510
rect 7012 37508 7036 37510
rect 7092 37508 7116 37510
rect 7172 37508 7196 37510
rect 7252 37508 7258 37510
rect 6950 37499 7258 37508
rect 11950 37564 12258 37573
rect 11950 37562 11956 37564
rect 12012 37562 12036 37564
rect 12092 37562 12116 37564
rect 12172 37562 12196 37564
rect 12252 37562 12258 37564
rect 12012 37510 12014 37562
rect 12194 37510 12196 37562
rect 11950 37508 11956 37510
rect 12012 37508 12036 37510
rect 12092 37508 12116 37510
rect 12172 37508 12196 37510
rect 12252 37508 12258 37510
rect 11950 37499 12258 37508
rect 16950 37564 17258 37573
rect 16950 37562 16956 37564
rect 17012 37562 17036 37564
rect 17092 37562 17116 37564
rect 17172 37562 17196 37564
rect 17252 37562 17258 37564
rect 17012 37510 17014 37562
rect 17194 37510 17196 37562
rect 16950 37508 16956 37510
rect 17012 37508 17036 37510
rect 17092 37508 17116 37510
rect 17172 37508 17196 37510
rect 17252 37508 17258 37510
rect 16950 37499 17258 37508
rect 21950 37564 22258 37573
rect 21950 37562 21956 37564
rect 22012 37562 22036 37564
rect 22092 37562 22116 37564
rect 22172 37562 22196 37564
rect 22252 37562 22258 37564
rect 22012 37510 22014 37562
rect 22194 37510 22196 37562
rect 21950 37508 21956 37510
rect 22012 37508 22036 37510
rect 22092 37508 22116 37510
rect 22172 37508 22196 37510
rect 22252 37508 22258 37510
rect 21950 37499 22258 37508
rect 26950 37564 27258 37573
rect 26950 37562 26956 37564
rect 27012 37562 27036 37564
rect 27092 37562 27116 37564
rect 27172 37562 27196 37564
rect 27252 37562 27258 37564
rect 27012 37510 27014 37562
rect 27194 37510 27196 37562
rect 26950 37508 26956 37510
rect 27012 37508 27036 37510
rect 27092 37508 27116 37510
rect 27172 37508 27196 37510
rect 27252 37508 27258 37510
rect 26950 37499 27258 37508
rect 31950 37564 32258 37573
rect 31950 37562 31956 37564
rect 32012 37562 32036 37564
rect 32092 37562 32116 37564
rect 32172 37562 32196 37564
rect 32252 37562 32258 37564
rect 32012 37510 32014 37562
rect 32194 37510 32196 37562
rect 31950 37508 31956 37510
rect 32012 37508 32036 37510
rect 32092 37508 32116 37510
rect 32172 37508 32196 37510
rect 32252 37508 32258 37510
rect 31950 37499 32258 37508
rect 36950 37564 37258 37573
rect 36950 37562 36956 37564
rect 37012 37562 37036 37564
rect 37092 37562 37116 37564
rect 37172 37562 37196 37564
rect 37252 37562 37258 37564
rect 37012 37510 37014 37562
rect 37194 37510 37196 37562
rect 36950 37508 36956 37510
rect 37012 37508 37036 37510
rect 37092 37508 37116 37510
rect 37172 37508 37196 37510
rect 37252 37508 37258 37510
rect 36950 37499 37258 37508
rect 2610 37020 2918 37029
rect 2610 37018 2616 37020
rect 2672 37018 2696 37020
rect 2752 37018 2776 37020
rect 2832 37018 2856 37020
rect 2912 37018 2918 37020
rect 2672 36966 2674 37018
rect 2854 36966 2856 37018
rect 2610 36964 2616 36966
rect 2672 36964 2696 36966
rect 2752 36964 2776 36966
rect 2832 36964 2856 36966
rect 2912 36964 2918 36966
rect 2610 36955 2918 36964
rect 7610 37020 7918 37029
rect 7610 37018 7616 37020
rect 7672 37018 7696 37020
rect 7752 37018 7776 37020
rect 7832 37018 7856 37020
rect 7912 37018 7918 37020
rect 7672 36966 7674 37018
rect 7854 36966 7856 37018
rect 7610 36964 7616 36966
rect 7672 36964 7696 36966
rect 7752 36964 7776 36966
rect 7832 36964 7856 36966
rect 7912 36964 7918 36966
rect 7610 36955 7918 36964
rect 12610 37020 12918 37029
rect 12610 37018 12616 37020
rect 12672 37018 12696 37020
rect 12752 37018 12776 37020
rect 12832 37018 12856 37020
rect 12912 37018 12918 37020
rect 12672 36966 12674 37018
rect 12854 36966 12856 37018
rect 12610 36964 12616 36966
rect 12672 36964 12696 36966
rect 12752 36964 12776 36966
rect 12832 36964 12856 36966
rect 12912 36964 12918 36966
rect 12610 36955 12918 36964
rect 17610 37020 17918 37029
rect 17610 37018 17616 37020
rect 17672 37018 17696 37020
rect 17752 37018 17776 37020
rect 17832 37018 17856 37020
rect 17912 37018 17918 37020
rect 17672 36966 17674 37018
rect 17854 36966 17856 37018
rect 17610 36964 17616 36966
rect 17672 36964 17696 36966
rect 17752 36964 17776 36966
rect 17832 36964 17856 36966
rect 17912 36964 17918 36966
rect 17610 36955 17918 36964
rect 22610 37020 22918 37029
rect 22610 37018 22616 37020
rect 22672 37018 22696 37020
rect 22752 37018 22776 37020
rect 22832 37018 22856 37020
rect 22912 37018 22918 37020
rect 22672 36966 22674 37018
rect 22854 36966 22856 37018
rect 22610 36964 22616 36966
rect 22672 36964 22696 36966
rect 22752 36964 22776 36966
rect 22832 36964 22856 36966
rect 22912 36964 22918 36966
rect 22610 36955 22918 36964
rect 27610 37020 27918 37029
rect 27610 37018 27616 37020
rect 27672 37018 27696 37020
rect 27752 37018 27776 37020
rect 27832 37018 27856 37020
rect 27912 37018 27918 37020
rect 27672 36966 27674 37018
rect 27854 36966 27856 37018
rect 27610 36964 27616 36966
rect 27672 36964 27696 36966
rect 27752 36964 27776 36966
rect 27832 36964 27856 36966
rect 27912 36964 27918 36966
rect 27610 36955 27918 36964
rect 32610 37020 32918 37029
rect 32610 37018 32616 37020
rect 32672 37018 32696 37020
rect 32752 37018 32776 37020
rect 32832 37018 32856 37020
rect 32912 37018 32918 37020
rect 32672 36966 32674 37018
rect 32854 36966 32856 37018
rect 32610 36964 32616 36966
rect 32672 36964 32696 36966
rect 32752 36964 32776 36966
rect 32832 36964 32856 36966
rect 32912 36964 32918 36966
rect 32610 36955 32918 36964
rect 37610 37020 37918 37029
rect 37610 37018 37616 37020
rect 37672 37018 37696 37020
rect 37752 37018 37776 37020
rect 37832 37018 37856 37020
rect 37912 37018 37918 37020
rect 37672 36966 37674 37018
rect 37854 36966 37856 37018
rect 37610 36964 37616 36966
rect 37672 36964 37696 36966
rect 37752 36964 37776 36966
rect 37832 36964 37856 36966
rect 37912 36964 37918 36966
rect 37610 36955 37918 36964
rect 1950 36476 2258 36485
rect 1950 36474 1956 36476
rect 2012 36474 2036 36476
rect 2092 36474 2116 36476
rect 2172 36474 2196 36476
rect 2252 36474 2258 36476
rect 2012 36422 2014 36474
rect 2194 36422 2196 36474
rect 1950 36420 1956 36422
rect 2012 36420 2036 36422
rect 2092 36420 2116 36422
rect 2172 36420 2196 36422
rect 2252 36420 2258 36422
rect 1950 36411 2258 36420
rect 6950 36476 7258 36485
rect 6950 36474 6956 36476
rect 7012 36474 7036 36476
rect 7092 36474 7116 36476
rect 7172 36474 7196 36476
rect 7252 36474 7258 36476
rect 7012 36422 7014 36474
rect 7194 36422 7196 36474
rect 6950 36420 6956 36422
rect 7012 36420 7036 36422
rect 7092 36420 7116 36422
rect 7172 36420 7196 36422
rect 7252 36420 7258 36422
rect 6950 36411 7258 36420
rect 11950 36476 12258 36485
rect 11950 36474 11956 36476
rect 12012 36474 12036 36476
rect 12092 36474 12116 36476
rect 12172 36474 12196 36476
rect 12252 36474 12258 36476
rect 12012 36422 12014 36474
rect 12194 36422 12196 36474
rect 11950 36420 11956 36422
rect 12012 36420 12036 36422
rect 12092 36420 12116 36422
rect 12172 36420 12196 36422
rect 12252 36420 12258 36422
rect 11950 36411 12258 36420
rect 16950 36476 17258 36485
rect 16950 36474 16956 36476
rect 17012 36474 17036 36476
rect 17092 36474 17116 36476
rect 17172 36474 17196 36476
rect 17252 36474 17258 36476
rect 17012 36422 17014 36474
rect 17194 36422 17196 36474
rect 16950 36420 16956 36422
rect 17012 36420 17036 36422
rect 17092 36420 17116 36422
rect 17172 36420 17196 36422
rect 17252 36420 17258 36422
rect 16950 36411 17258 36420
rect 21950 36476 22258 36485
rect 21950 36474 21956 36476
rect 22012 36474 22036 36476
rect 22092 36474 22116 36476
rect 22172 36474 22196 36476
rect 22252 36474 22258 36476
rect 22012 36422 22014 36474
rect 22194 36422 22196 36474
rect 21950 36420 21956 36422
rect 22012 36420 22036 36422
rect 22092 36420 22116 36422
rect 22172 36420 22196 36422
rect 22252 36420 22258 36422
rect 21950 36411 22258 36420
rect 26950 36476 27258 36485
rect 26950 36474 26956 36476
rect 27012 36474 27036 36476
rect 27092 36474 27116 36476
rect 27172 36474 27196 36476
rect 27252 36474 27258 36476
rect 27012 36422 27014 36474
rect 27194 36422 27196 36474
rect 26950 36420 26956 36422
rect 27012 36420 27036 36422
rect 27092 36420 27116 36422
rect 27172 36420 27196 36422
rect 27252 36420 27258 36422
rect 26950 36411 27258 36420
rect 31950 36476 32258 36485
rect 31950 36474 31956 36476
rect 32012 36474 32036 36476
rect 32092 36474 32116 36476
rect 32172 36474 32196 36476
rect 32252 36474 32258 36476
rect 32012 36422 32014 36474
rect 32194 36422 32196 36474
rect 31950 36420 31956 36422
rect 32012 36420 32036 36422
rect 32092 36420 32116 36422
rect 32172 36420 32196 36422
rect 32252 36420 32258 36422
rect 31950 36411 32258 36420
rect 36950 36476 37258 36485
rect 36950 36474 36956 36476
rect 37012 36474 37036 36476
rect 37092 36474 37116 36476
rect 37172 36474 37196 36476
rect 37252 36474 37258 36476
rect 37012 36422 37014 36474
rect 37194 36422 37196 36474
rect 36950 36420 36956 36422
rect 37012 36420 37036 36422
rect 37092 36420 37116 36422
rect 37172 36420 37196 36422
rect 37252 36420 37258 36422
rect 36950 36411 37258 36420
rect 2610 35932 2918 35941
rect 2610 35930 2616 35932
rect 2672 35930 2696 35932
rect 2752 35930 2776 35932
rect 2832 35930 2856 35932
rect 2912 35930 2918 35932
rect 2672 35878 2674 35930
rect 2854 35878 2856 35930
rect 2610 35876 2616 35878
rect 2672 35876 2696 35878
rect 2752 35876 2776 35878
rect 2832 35876 2856 35878
rect 2912 35876 2918 35878
rect 2610 35867 2918 35876
rect 7610 35932 7918 35941
rect 7610 35930 7616 35932
rect 7672 35930 7696 35932
rect 7752 35930 7776 35932
rect 7832 35930 7856 35932
rect 7912 35930 7918 35932
rect 7672 35878 7674 35930
rect 7854 35878 7856 35930
rect 7610 35876 7616 35878
rect 7672 35876 7696 35878
rect 7752 35876 7776 35878
rect 7832 35876 7856 35878
rect 7912 35876 7918 35878
rect 7610 35867 7918 35876
rect 12610 35932 12918 35941
rect 12610 35930 12616 35932
rect 12672 35930 12696 35932
rect 12752 35930 12776 35932
rect 12832 35930 12856 35932
rect 12912 35930 12918 35932
rect 12672 35878 12674 35930
rect 12854 35878 12856 35930
rect 12610 35876 12616 35878
rect 12672 35876 12696 35878
rect 12752 35876 12776 35878
rect 12832 35876 12856 35878
rect 12912 35876 12918 35878
rect 12610 35867 12918 35876
rect 17610 35932 17918 35941
rect 17610 35930 17616 35932
rect 17672 35930 17696 35932
rect 17752 35930 17776 35932
rect 17832 35930 17856 35932
rect 17912 35930 17918 35932
rect 17672 35878 17674 35930
rect 17854 35878 17856 35930
rect 17610 35876 17616 35878
rect 17672 35876 17696 35878
rect 17752 35876 17776 35878
rect 17832 35876 17856 35878
rect 17912 35876 17918 35878
rect 17610 35867 17918 35876
rect 22610 35932 22918 35941
rect 22610 35930 22616 35932
rect 22672 35930 22696 35932
rect 22752 35930 22776 35932
rect 22832 35930 22856 35932
rect 22912 35930 22918 35932
rect 22672 35878 22674 35930
rect 22854 35878 22856 35930
rect 22610 35876 22616 35878
rect 22672 35876 22696 35878
rect 22752 35876 22776 35878
rect 22832 35876 22856 35878
rect 22912 35876 22918 35878
rect 22610 35867 22918 35876
rect 27610 35932 27918 35941
rect 27610 35930 27616 35932
rect 27672 35930 27696 35932
rect 27752 35930 27776 35932
rect 27832 35930 27856 35932
rect 27912 35930 27918 35932
rect 27672 35878 27674 35930
rect 27854 35878 27856 35930
rect 27610 35876 27616 35878
rect 27672 35876 27696 35878
rect 27752 35876 27776 35878
rect 27832 35876 27856 35878
rect 27912 35876 27918 35878
rect 27610 35867 27918 35876
rect 32610 35932 32918 35941
rect 32610 35930 32616 35932
rect 32672 35930 32696 35932
rect 32752 35930 32776 35932
rect 32832 35930 32856 35932
rect 32912 35930 32918 35932
rect 32672 35878 32674 35930
rect 32854 35878 32856 35930
rect 32610 35876 32616 35878
rect 32672 35876 32696 35878
rect 32752 35876 32776 35878
rect 32832 35876 32856 35878
rect 32912 35876 32918 35878
rect 32610 35867 32918 35876
rect 37610 35932 37918 35941
rect 37610 35930 37616 35932
rect 37672 35930 37696 35932
rect 37752 35930 37776 35932
rect 37832 35930 37856 35932
rect 37912 35930 37918 35932
rect 37672 35878 37674 35930
rect 37854 35878 37856 35930
rect 37610 35876 37616 35878
rect 37672 35876 37696 35878
rect 37752 35876 37776 35878
rect 37832 35876 37856 35878
rect 37912 35876 37918 35878
rect 37610 35867 37918 35876
rect 1950 35388 2258 35397
rect 1950 35386 1956 35388
rect 2012 35386 2036 35388
rect 2092 35386 2116 35388
rect 2172 35386 2196 35388
rect 2252 35386 2258 35388
rect 2012 35334 2014 35386
rect 2194 35334 2196 35386
rect 1950 35332 1956 35334
rect 2012 35332 2036 35334
rect 2092 35332 2116 35334
rect 2172 35332 2196 35334
rect 2252 35332 2258 35334
rect 1950 35323 2258 35332
rect 6950 35388 7258 35397
rect 6950 35386 6956 35388
rect 7012 35386 7036 35388
rect 7092 35386 7116 35388
rect 7172 35386 7196 35388
rect 7252 35386 7258 35388
rect 7012 35334 7014 35386
rect 7194 35334 7196 35386
rect 6950 35332 6956 35334
rect 7012 35332 7036 35334
rect 7092 35332 7116 35334
rect 7172 35332 7196 35334
rect 7252 35332 7258 35334
rect 6950 35323 7258 35332
rect 11950 35388 12258 35397
rect 11950 35386 11956 35388
rect 12012 35386 12036 35388
rect 12092 35386 12116 35388
rect 12172 35386 12196 35388
rect 12252 35386 12258 35388
rect 12012 35334 12014 35386
rect 12194 35334 12196 35386
rect 11950 35332 11956 35334
rect 12012 35332 12036 35334
rect 12092 35332 12116 35334
rect 12172 35332 12196 35334
rect 12252 35332 12258 35334
rect 11950 35323 12258 35332
rect 16950 35388 17258 35397
rect 16950 35386 16956 35388
rect 17012 35386 17036 35388
rect 17092 35386 17116 35388
rect 17172 35386 17196 35388
rect 17252 35386 17258 35388
rect 17012 35334 17014 35386
rect 17194 35334 17196 35386
rect 16950 35332 16956 35334
rect 17012 35332 17036 35334
rect 17092 35332 17116 35334
rect 17172 35332 17196 35334
rect 17252 35332 17258 35334
rect 16950 35323 17258 35332
rect 21950 35388 22258 35397
rect 21950 35386 21956 35388
rect 22012 35386 22036 35388
rect 22092 35386 22116 35388
rect 22172 35386 22196 35388
rect 22252 35386 22258 35388
rect 22012 35334 22014 35386
rect 22194 35334 22196 35386
rect 21950 35332 21956 35334
rect 22012 35332 22036 35334
rect 22092 35332 22116 35334
rect 22172 35332 22196 35334
rect 22252 35332 22258 35334
rect 21950 35323 22258 35332
rect 26950 35388 27258 35397
rect 26950 35386 26956 35388
rect 27012 35386 27036 35388
rect 27092 35386 27116 35388
rect 27172 35386 27196 35388
rect 27252 35386 27258 35388
rect 27012 35334 27014 35386
rect 27194 35334 27196 35386
rect 26950 35332 26956 35334
rect 27012 35332 27036 35334
rect 27092 35332 27116 35334
rect 27172 35332 27196 35334
rect 27252 35332 27258 35334
rect 26950 35323 27258 35332
rect 31950 35388 32258 35397
rect 31950 35386 31956 35388
rect 32012 35386 32036 35388
rect 32092 35386 32116 35388
rect 32172 35386 32196 35388
rect 32252 35386 32258 35388
rect 32012 35334 32014 35386
rect 32194 35334 32196 35386
rect 31950 35332 31956 35334
rect 32012 35332 32036 35334
rect 32092 35332 32116 35334
rect 32172 35332 32196 35334
rect 32252 35332 32258 35334
rect 31950 35323 32258 35332
rect 36950 35388 37258 35397
rect 36950 35386 36956 35388
rect 37012 35386 37036 35388
rect 37092 35386 37116 35388
rect 37172 35386 37196 35388
rect 37252 35386 37258 35388
rect 37012 35334 37014 35386
rect 37194 35334 37196 35386
rect 36950 35332 36956 35334
rect 37012 35332 37036 35334
rect 37092 35332 37116 35334
rect 37172 35332 37196 35334
rect 37252 35332 37258 35334
rect 36950 35323 37258 35332
rect 2610 34844 2918 34853
rect 2610 34842 2616 34844
rect 2672 34842 2696 34844
rect 2752 34842 2776 34844
rect 2832 34842 2856 34844
rect 2912 34842 2918 34844
rect 2672 34790 2674 34842
rect 2854 34790 2856 34842
rect 2610 34788 2616 34790
rect 2672 34788 2696 34790
rect 2752 34788 2776 34790
rect 2832 34788 2856 34790
rect 2912 34788 2918 34790
rect 2610 34779 2918 34788
rect 7610 34844 7918 34853
rect 7610 34842 7616 34844
rect 7672 34842 7696 34844
rect 7752 34842 7776 34844
rect 7832 34842 7856 34844
rect 7912 34842 7918 34844
rect 7672 34790 7674 34842
rect 7854 34790 7856 34842
rect 7610 34788 7616 34790
rect 7672 34788 7696 34790
rect 7752 34788 7776 34790
rect 7832 34788 7856 34790
rect 7912 34788 7918 34790
rect 7610 34779 7918 34788
rect 12610 34844 12918 34853
rect 12610 34842 12616 34844
rect 12672 34842 12696 34844
rect 12752 34842 12776 34844
rect 12832 34842 12856 34844
rect 12912 34842 12918 34844
rect 12672 34790 12674 34842
rect 12854 34790 12856 34842
rect 12610 34788 12616 34790
rect 12672 34788 12696 34790
rect 12752 34788 12776 34790
rect 12832 34788 12856 34790
rect 12912 34788 12918 34790
rect 12610 34779 12918 34788
rect 17610 34844 17918 34853
rect 17610 34842 17616 34844
rect 17672 34842 17696 34844
rect 17752 34842 17776 34844
rect 17832 34842 17856 34844
rect 17912 34842 17918 34844
rect 17672 34790 17674 34842
rect 17854 34790 17856 34842
rect 17610 34788 17616 34790
rect 17672 34788 17696 34790
rect 17752 34788 17776 34790
rect 17832 34788 17856 34790
rect 17912 34788 17918 34790
rect 17610 34779 17918 34788
rect 22610 34844 22918 34853
rect 22610 34842 22616 34844
rect 22672 34842 22696 34844
rect 22752 34842 22776 34844
rect 22832 34842 22856 34844
rect 22912 34842 22918 34844
rect 22672 34790 22674 34842
rect 22854 34790 22856 34842
rect 22610 34788 22616 34790
rect 22672 34788 22696 34790
rect 22752 34788 22776 34790
rect 22832 34788 22856 34790
rect 22912 34788 22918 34790
rect 22610 34779 22918 34788
rect 27610 34844 27918 34853
rect 27610 34842 27616 34844
rect 27672 34842 27696 34844
rect 27752 34842 27776 34844
rect 27832 34842 27856 34844
rect 27912 34842 27918 34844
rect 27672 34790 27674 34842
rect 27854 34790 27856 34842
rect 27610 34788 27616 34790
rect 27672 34788 27696 34790
rect 27752 34788 27776 34790
rect 27832 34788 27856 34790
rect 27912 34788 27918 34790
rect 27610 34779 27918 34788
rect 32610 34844 32918 34853
rect 32610 34842 32616 34844
rect 32672 34842 32696 34844
rect 32752 34842 32776 34844
rect 32832 34842 32856 34844
rect 32912 34842 32918 34844
rect 32672 34790 32674 34842
rect 32854 34790 32856 34842
rect 32610 34788 32616 34790
rect 32672 34788 32696 34790
rect 32752 34788 32776 34790
rect 32832 34788 32856 34790
rect 32912 34788 32918 34790
rect 32610 34779 32918 34788
rect 37610 34844 37918 34853
rect 37610 34842 37616 34844
rect 37672 34842 37696 34844
rect 37752 34842 37776 34844
rect 37832 34842 37856 34844
rect 37912 34842 37918 34844
rect 37672 34790 37674 34842
rect 37854 34790 37856 34842
rect 37610 34788 37616 34790
rect 37672 34788 37696 34790
rect 37752 34788 37776 34790
rect 37832 34788 37856 34790
rect 37912 34788 37918 34790
rect 37610 34779 37918 34788
rect 1950 34300 2258 34309
rect 1950 34298 1956 34300
rect 2012 34298 2036 34300
rect 2092 34298 2116 34300
rect 2172 34298 2196 34300
rect 2252 34298 2258 34300
rect 2012 34246 2014 34298
rect 2194 34246 2196 34298
rect 1950 34244 1956 34246
rect 2012 34244 2036 34246
rect 2092 34244 2116 34246
rect 2172 34244 2196 34246
rect 2252 34244 2258 34246
rect 1950 34235 2258 34244
rect 6950 34300 7258 34309
rect 6950 34298 6956 34300
rect 7012 34298 7036 34300
rect 7092 34298 7116 34300
rect 7172 34298 7196 34300
rect 7252 34298 7258 34300
rect 7012 34246 7014 34298
rect 7194 34246 7196 34298
rect 6950 34244 6956 34246
rect 7012 34244 7036 34246
rect 7092 34244 7116 34246
rect 7172 34244 7196 34246
rect 7252 34244 7258 34246
rect 6950 34235 7258 34244
rect 11950 34300 12258 34309
rect 11950 34298 11956 34300
rect 12012 34298 12036 34300
rect 12092 34298 12116 34300
rect 12172 34298 12196 34300
rect 12252 34298 12258 34300
rect 12012 34246 12014 34298
rect 12194 34246 12196 34298
rect 11950 34244 11956 34246
rect 12012 34244 12036 34246
rect 12092 34244 12116 34246
rect 12172 34244 12196 34246
rect 12252 34244 12258 34246
rect 11950 34235 12258 34244
rect 16950 34300 17258 34309
rect 16950 34298 16956 34300
rect 17012 34298 17036 34300
rect 17092 34298 17116 34300
rect 17172 34298 17196 34300
rect 17252 34298 17258 34300
rect 17012 34246 17014 34298
rect 17194 34246 17196 34298
rect 16950 34244 16956 34246
rect 17012 34244 17036 34246
rect 17092 34244 17116 34246
rect 17172 34244 17196 34246
rect 17252 34244 17258 34246
rect 16950 34235 17258 34244
rect 21950 34300 22258 34309
rect 21950 34298 21956 34300
rect 22012 34298 22036 34300
rect 22092 34298 22116 34300
rect 22172 34298 22196 34300
rect 22252 34298 22258 34300
rect 22012 34246 22014 34298
rect 22194 34246 22196 34298
rect 21950 34244 21956 34246
rect 22012 34244 22036 34246
rect 22092 34244 22116 34246
rect 22172 34244 22196 34246
rect 22252 34244 22258 34246
rect 21950 34235 22258 34244
rect 26950 34300 27258 34309
rect 26950 34298 26956 34300
rect 27012 34298 27036 34300
rect 27092 34298 27116 34300
rect 27172 34298 27196 34300
rect 27252 34298 27258 34300
rect 27012 34246 27014 34298
rect 27194 34246 27196 34298
rect 26950 34244 26956 34246
rect 27012 34244 27036 34246
rect 27092 34244 27116 34246
rect 27172 34244 27196 34246
rect 27252 34244 27258 34246
rect 26950 34235 27258 34244
rect 31950 34300 32258 34309
rect 31950 34298 31956 34300
rect 32012 34298 32036 34300
rect 32092 34298 32116 34300
rect 32172 34298 32196 34300
rect 32252 34298 32258 34300
rect 32012 34246 32014 34298
rect 32194 34246 32196 34298
rect 31950 34244 31956 34246
rect 32012 34244 32036 34246
rect 32092 34244 32116 34246
rect 32172 34244 32196 34246
rect 32252 34244 32258 34246
rect 31950 34235 32258 34244
rect 36950 34300 37258 34309
rect 36950 34298 36956 34300
rect 37012 34298 37036 34300
rect 37092 34298 37116 34300
rect 37172 34298 37196 34300
rect 37252 34298 37258 34300
rect 37012 34246 37014 34298
rect 37194 34246 37196 34298
rect 36950 34244 36956 34246
rect 37012 34244 37036 34246
rect 37092 34244 37116 34246
rect 37172 34244 37196 34246
rect 37252 34244 37258 34246
rect 36950 34235 37258 34244
rect 2610 33756 2918 33765
rect 2610 33754 2616 33756
rect 2672 33754 2696 33756
rect 2752 33754 2776 33756
rect 2832 33754 2856 33756
rect 2912 33754 2918 33756
rect 2672 33702 2674 33754
rect 2854 33702 2856 33754
rect 2610 33700 2616 33702
rect 2672 33700 2696 33702
rect 2752 33700 2776 33702
rect 2832 33700 2856 33702
rect 2912 33700 2918 33702
rect 2610 33691 2918 33700
rect 7610 33756 7918 33765
rect 7610 33754 7616 33756
rect 7672 33754 7696 33756
rect 7752 33754 7776 33756
rect 7832 33754 7856 33756
rect 7912 33754 7918 33756
rect 7672 33702 7674 33754
rect 7854 33702 7856 33754
rect 7610 33700 7616 33702
rect 7672 33700 7696 33702
rect 7752 33700 7776 33702
rect 7832 33700 7856 33702
rect 7912 33700 7918 33702
rect 7610 33691 7918 33700
rect 12610 33756 12918 33765
rect 12610 33754 12616 33756
rect 12672 33754 12696 33756
rect 12752 33754 12776 33756
rect 12832 33754 12856 33756
rect 12912 33754 12918 33756
rect 12672 33702 12674 33754
rect 12854 33702 12856 33754
rect 12610 33700 12616 33702
rect 12672 33700 12696 33702
rect 12752 33700 12776 33702
rect 12832 33700 12856 33702
rect 12912 33700 12918 33702
rect 12610 33691 12918 33700
rect 17610 33756 17918 33765
rect 17610 33754 17616 33756
rect 17672 33754 17696 33756
rect 17752 33754 17776 33756
rect 17832 33754 17856 33756
rect 17912 33754 17918 33756
rect 17672 33702 17674 33754
rect 17854 33702 17856 33754
rect 17610 33700 17616 33702
rect 17672 33700 17696 33702
rect 17752 33700 17776 33702
rect 17832 33700 17856 33702
rect 17912 33700 17918 33702
rect 17610 33691 17918 33700
rect 22610 33756 22918 33765
rect 22610 33754 22616 33756
rect 22672 33754 22696 33756
rect 22752 33754 22776 33756
rect 22832 33754 22856 33756
rect 22912 33754 22918 33756
rect 22672 33702 22674 33754
rect 22854 33702 22856 33754
rect 22610 33700 22616 33702
rect 22672 33700 22696 33702
rect 22752 33700 22776 33702
rect 22832 33700 22856 33702
rect 22912 33700 22918 33702
rect 22610 33691 22918 33700
rect 27610 33756 27918 33765
rect 27610 33754 27616 33756
rect 27672 33754 27696 33756
rect 27752 33754 27776 33756
rect 27832 33754 27856 33756
rect 27912 33754 27918 33756
rect 27672 33702 27674 33754
rect 27854 33702 27856 33754
rect 27610 33700 27616 33702
rect 27672 33700 27696 33702
rect 27752 33700 27776 33702
rect 27832 33700 27856 33702
rect 27912 33700 27918 33702
rect 27610 33691 27918 33700
rect 32610 33756 32918 33765
rect 32610 33754 32616 33756
rect 32672 33754 32696 33756
rect 32752 33754 32776 33756
rect 32832 33754 32856 33756
rect 32912 33754 32918 33756
rect 32672 33702 32674 33754
rect 32854 33702 32856 33754
rect 32610 33700 32616 33702
rect 32672 33700 32696 33702
rect 32752 33700 32776 33702
rect 32832 33700 32856 33702
rect 32912 33700 32918 33702
rect 32610 33691 32918 33700
rect 37610 33756 37918 33765
rect 37610 33754 37616 33756
rect 37672 33754 37696 33756
rect 37752 33754 37776 33756
rect 37832 33754 37856 33756
rect 37912 33754 37918 33756
rect 37672 33702 37674 33754
rect 37854 33702 37856 33754
rect 37610 33700 37616 33702
rect 37672 33700 37696 33702
rect 37752 33700 37776 33702
rect 37832 33700 37856 33702
rect 37912 33700 37918 33702
rect 37610 33691 37918 33700
rect 1950 33212 2258 33221
rect 1950 33210 1956 33212
rect 2012 33210 2036 33212
rect 2092 33210 2116 33212
rect 2172 33210 2196 33212
rect 2252 33210 2258 33212
rect 2012 33158 2014 33210
rect 2194 33158 2196 33210
rect 1950 33156 1956 33158
rect 2012 33156 2036 33158
rect 2092 33156 2116 33158
rect 2172 33156 2196 33158
rect 2252 33156 2258 33158
rect 1950 33147 2258 33156
rect 6950 33212 7258 33221
rect 6950 33210 6956 33212
rect 7012 33210 7036 33212
rect 7092 33210 7116 33212
rect 7172 33210 7196 33212
rect 7252 33210 7258 33212
rect 7012 33158 7014 33210
rect 7194 33158 7196 33210
rect 6950 33156 6956 33158
rect 7012 33156 7036 33158
rect 7092 33156 7116 33158
rect 7172 33156 7196 33158
rect 7252 33156 7258 33158
rect 6950 33147 7258 33156
rect 11950 33212 12258 33221
rect 11950 33210 11956 33212
rect 12012 33210 12036 33212
rect 12092 33210 12116 33212
rect 12172 33210 12196 33212
rect 12252 33210 12258 33212
rect 12012 33158 12014 33210
rect 12194 33158 12196 33210
rect 11950 33156 11956 33158
rect 12012 33156 12036 33158
rect 12092 33156 12116 33158
rect 12172 33156 12196 33158
rect 12252 33156 12258 33158
rect 11950 33147 12258 33156
rect 16950 33212 17258 33221
rect 16950 33210 16956 33212
rect 17012 33210 17036 33212
rect 17092 33210 17116 33212
rect 17172 33210 17196 33212
rect 17252 33210 17258 33212
rect 17012 33158 17014 33210
rect 17194 33158 17196 33210
rect 16950 33156 16956 33158
rect 17012 33156 17036 33158
rect 17092 33156 17116 33158
rect 17172 33156 17196 33158
rect 17252 33156 17258 33158
rect 16950 33147 17258 33156
rect 21950 33212 22258 33221
rect 21950 33210 21956 33212
rect 22012 33210 22036 33212
rect 22092 33210 22116 33212
rect 22172 33210 22196 33212
rect 22252 33210 22258 33212
rect 22012 33158 22014 33210
rect 22194 33158 22196 33210
rect 21950 33156 21956 33158
rect 22012 33156 22036 33158
rect 22092 33156 22116 33158
rect 22172 33156 22196 33158
rect 22252 33156 22258 33158
rect 21950 33147 22258 33156
rect 26950 33212 27258 33221
rect 26950 33210 26956 33212
rect 27012 33210 27036 33212
rect 27092 33210 27116 33212
rect 27172 33210 27196 33212
rect 27252 33210 27258 33212
rect 27012 33158 27014 33210
rect 27194 33158 27196 33210
rect 26950 33156 26956 33158
rect 27012 33156 27036 33158
rect 27092 33156 27116 33158
rect 27172 33156 27196 33158
rect 27252 33156 27258 33158
rect 26950 33147 27258 33156
rect 31950 33212 32258 33221
rect 31950 33210 31956 33212
rect 32012 33210 32036 33212
rect 32092 33210 32116 33212
rect 32172 33210 32196 33212
rect 32252 33210 32258 33212
rect 32012 33158 32014 33210
rect 32194 33158 32196 33210
rect 31950 33156 31956 33158
rect 32012 33156 32036 33158
rect 32092 33156 32116 33158
rect 32172 33156 32196 33158
rect 32252 33156 32258 33158
rect 31950 33147 32258 33156
rect 36950 33212 37258 33221
rect 36950 33210 36956 33212
rect 37012 33210 37036 33212
rect 37092 33210 37116 33212
rect 37172 33210 37196 33212
rect 37252 33210 37258 33212
rect 37012 33158 37014 33210
rect 37194 33158 37196 33210
rect 36950 33156 36956 33158
rect 37012 33156 37036 33158
rect 37092 33156 37116 33158
rect 37172 33156 37196 33158
rect 37252 33156 37258 33158
rect 36950 33147 37258 33156
rect 2610 32668 2918 32677
rect 2610 32666 2616 32668
rect 2672 32666 2696 32668
rect 2752 32666 2776 32668
rect 2832 32666 2856 32668
rect 2912 32666 2918 32668
rect 2672 32614 2674 32666
rect 2854 32614 2856 32666
rect 2610 32612 2616 32614
rect 2672 32612 2696 32614
rect 2752 32612 2776 32614
rect 2832 32612 2856 32614
rect 2912 32612 2918 32614
rect 2610 32603 2918 32612
rect 7610 32668 7918 32677
rect 7610 32666 7616 32668
rect 7672 32666 7696 32668
rect 7752 32666 7776 32668
rect 7832 32666 7856 32668
rect 7912 32666 7918 32668
rect 7672 32614 7674 32666
rect 7854 32614 7856 32666
rect 7610 32612 7616 32614
rect 7672 32612 7696 32614
rect 7752 32612 7776 32614
rect 7832 32612 7856 32614
rect 7912 32612 7918 32614
rect 7610 32603 7918 32612
rect 12610 32668 12918 32677
rect 12610 32666 12616 32668
rect 12672 32666 12696 32668
rect 12752 32666 12776 32668
rect 12832 32666 12856 32668
rect 12912 32666 12918 32668
rect 12672 32614 12674 32666
rect 12854 32614 12856 32666
rect 12610 32612 12616 32614
rect 12672 32612 12696 32614
rect 12752 32612 12776 32614
rect 12832 32612 12856 32614
rect 12912 32612 12918 32614
rect 12610 32603 12918 32612
rect 17610 32668 17918 32677
rect 17610 32666 17616 32668
rect 17672 32666 17696 32668
rect 17752 32666 17776 32668
rect 17832 32666 17856 32668
rect 17912 32666 17918 32668
rect 17672 32614 17674 32666
rect 17854 32614 17856 32666
rect 17610 32612 17616 32614
rect 17672 32612 17696 32614
rect 17752 32612 17776 32614
rect 17832 32612 17856 32614
rect 17912 32612 17918 32614
rect 17610 32603 17918 32612
rect 22610 32668 22918 32677
rect 22610 32666 22616 32668
rect 22672 32666 22696 32668
rect 22752 32666 22776 32668
rect 22832 32666 22856 32668
rect 22912 32666 22918 32668
rect 22672 32614 22674 32666
rect 22854 32614 22856 32666
rect 22610 32612 22616 32614
rect 22672 32612 22696 32614
rect 22752 32612 22776 32614
rect 22832 32612 22856 32614
rect 22912 32612 22918 32614
rect 22610 32603 22918 32612
rect 27610 32668 27918 32677
rect 27610 32666 27616 32668
rect 27672 32666 27696 32668
rect 27752 32666 27776 32668
rect 27832 32666 27856 32668
rect 27912 32666 27918 32668
rect 27672 32614 27674 32666
rect 27854 32614 27856 32666
rect 27610 32612 27616 32614
rect 27672 32612 27696 32614
rect 27752 32612 27776 32614
rect 27832 32612 27856 32614
rect 27912 32612 27918 32614
rect 27610 32603 27918 32612
rect 32610 32668 32918 32677
rect 32610 32666 32616 32668
rect 32672 32666 32696 32668
rect 32752 32666 32776 32668
rect 32832 32666 32856 32668
rect 32912 32666 32918 32668
rect 32672 32614 32674 32666
rect 32854 32614 32856 32666
rect 32610 32612 32616 32614
rect 32672 32612 32696 32614
rect 32752 32612 32776 32614
rect 32832 32612 32856 32614
rect 32912 32612 32918 32614
rect 32610 32603 32918 32612
rect 37610 32668 37918 32677
rect 37610 32666 37616 32668
rect 37672 32666 37696 32668
rect 37752 32666 37776 32668
rect 37832 32666 37856 32668
rect 37912 32666 37918 32668
rect 37672 32614 37674 32666
rect 37854 32614 37856 32666
rect 37610 32612 37616 32614
rect 37672 32612 37696 32614
rect 37752 32612 37776 32614
rect 37832 32612 37856 32614
rect 37912 32612 37918 32614
rect 37610 32603 37918 32612
rect 1950 32124 2258 32133
rect 1950 32122 1956 32124
rect 2012 32122 2036 32124
rect 2092 32122 2116 32124
rect 2172 32122 2196 32124
rect 2252 32122 2258 32124
rect 2012 32070 2014 32122
rect 2194 32070 2196 32122
rect 1950 32068 1956 32070
rect 2012 32068 2036 32070
rect 2092 32068 2116 32070
rect 2172 32068 2196 32070
rect 2252 32068 2258 32070
rect 1950 32059 2258 32068
rect 6950 32124 7258 32133
rect 6950 32122 6956 32124
rect 7012 32122 7036 32124
rect 7092 32122 7116 32124
rect 7172 32122 7196 32124
rect 7252 32122 7258 32124
rect 7012 32070 7014 32122
rect 7194 32070 7196 32122
rect 6950 32068 6956 32070
rect 7012 32068 7036 32070
rect 7092 32068 7116 32070
rect 7172 32068 7196 32070
rect 7252 32068 7258 32070
rect 6950 32059 7258 32068
rect 11950 32124 12258 32133
rect 11950 32122 11956 32124
rect 12012 32122 12036 32124
rect 12092 32122 12116 32124
rect 12172 32122 12196 32124
rect 12252 32122 12258 32124
rect 12012 32070 12014 32122
rect 12194 32070 12196 32122
rect 11950 32068 11956 32070
rect 12012 32068 12036 32070
rect 12092 32068 12116 32070
rect 12172 32068 12196 32070
rect 12252 32068 12258 32070
rect 11950 32059 12258 32068
rect 16950 32124 17258 32133
rect 16950 32122 16956 32124
rect 17012 32122 17036 32124
rect 17092 32122 17116 32124
rect 17172 32122 17196 32124
rect 17252 32122 17258 32124
rect 17012 32070 17014 32122
rect 17194 32070 17196 32122
rect 16950 32068 16956 32070
rect 17012 32068 17036 32070
rect 17092 32068 17116 32070
rect 17172 32068 17196 32070
rect 17252 32068 17258 32070
rect 16950 32059 17258 32068
rect 21950 32124 22258 32133
rect 21950 32122 21956 32124
rect 22012 32122 22036 32124
rect 22092 32122 22116 32124
rect 22172 32122 22196 32124
rect 22252 32122 22258 32124
rect 22012 32070 22014 32122
rect 22194 32070 22196 32122
rect 21950 32068 21956 32070
rect 22012 32068 22036 32070
rect 22092 32068 22116 32070
rect 22172 32068 22196 32070
rect 22252 32068 22258 32070
rect 21950 32059 22258 32068
rect 26950 32124 27258 32133
rect 26950 32122 26956 32124
rect 27012 32122 27036 32124
rect 27092 32122 27116 32124
rect 27172 32122 27196 32124
rect 27252 32122 27258 32124
rect 27012 32070 27014 32122
rect 27194 32070 27196 32122
rect 26950 32068 26956 32070
rect 27012 32068 27036 32070
rect 27092 32068 27116 32070
rect 27172 32068 27196 32070
rect 27252 32068 27258 32070
rect 26950 32059 27258 32068
rect 31950 32124 32258 32133
rect 31950 32122 31956 32124
rect 32012 32122 32036 32124
rect 32092 32122 32116 32124
rect 32172 32122 32196 32124
rect 32252 32122 32258 32124
rect 32012 32070 32014 32122
rect 32194 32070 32196 32122
rect 31950 32068 31956 32070
rect 32012 32068 32036 32070
rect 32092 32068 32116 32070
rect 32172 32068 32196 32070
rect 32252 32068 32258 32070
rect 31950 32059 32258 32068
rect 36950 32124 37258 32133
rect 36950 32122 36956 32124
rect 37012 32122 37036 32124
rect 37092 32122 37116 32124
rect 37172 32122 37196 32124
rect 37252 32122 37258 32124
rect 37012 32070 37014 32122
rect 37194 32070 37196 32122
rect 36950 32068 36956 32070
rect 37012 32068 37036 32070
rect 37092 32068 37116 32070
rect 37172 32068 37196 32070
rect 37252 32068 37258 32070
rect 36950 32059 37258 32068
rect 2610 31580 2918 31589
rect 2610 31578 2616 31580
rect 2672 31578 2696 31580
rect 2752 31578 2776 31580
rect 2832 31578 2856 31580
rect 2912 31578 2918 31580
rect 2672 31526 2674 31578
rect 2854 31526 2856 31578
rect 2610 31524 2616 31526
rect 2672 31524 2696 31526
rect 2752 31524 2776 31526
rect 2832 31524 2856 31526
rect 2912 31524 2918 31526
rect 2610 31515 2918 31524
rect 7610 31580 7918 31589
rect 7610 31578 7616 31580
rect 7672 31578 7696 31580
rect 7752 31578 7776 31580
rect 7832 31578 7856 31580
rect 7912 31578 7918 31580
rect 7672 31526 7674 31578
rect 7854 31526 7856 31578
rect 7610 31524 7616 31526
rect 7672 31524 7696 31526
rect 7752 31524 7776 31526
rect 7832 31524 7856 31526
rect 7912 31524 7918 31526
rect 7610 31515 7918 31524
rect 12610 31580 12918 31589
rect 12610 31578 12616 31580
rect 12672 31578 12696 31580
rect 12752 31578 12776 31580
rect 12832 31578 12856 31580
rect 12912 31578 12918 31580
rect 12672 31526 12674 31578
rect 12854 31526 12856 31578
rect 12610 31524 12616 31526
rect 12672 31524 12696 31526
rect 12752 31524 12776 31526
rect 12832 31524 12856 31526
rect 12912 31524 12918 31526
rect 12610 31515 12918 31524
rect 17610 31580 17918 31589
rect 17610 31578 17616 31580
rect 17672 31578 17696 31580
rect 17752 31578 17776 31580
rect 17832 31578 17856 31580
rect 17912 31578 17918 31580
rect 17672 31526 17674 31578
rect 17854 31526 17856 31578
rect 17610 31524 17616 31526
rect 17672 31524 17696 31526
rect 17752 31524 17776 31526
rect 17832 31524 17856 31526
rect 17912 31524 17918 31526
rect 17610 31515 17918 31524
rect 22610 31580 22918 31589
rect 22610 31578 22616 31580
rect 22672 31578 22696 31580
rect 22752 31578 22776 31580
rect 22832 31578 22856 31580
rect 22912 31578 22918 31580
rect 22672 31526 22674 31578
rect 22854 31526 22856 31578
rect 22610 31524 22616 31526
rect 22672 31524 22696 31526
rect 22752 31524 22776 31526
rect 22832 31524 22856 31526
rect 22912 31524 22918 31526
rect 22610 31515 22918 31524
rect 27610 31580 27918 31589
rect 27610 31578 27616 31580
rect 27672 31578 27696 31580
rect 27752 31578 27776 31580
rect 27832 31578 27856 31580
rect 27912 31578 27918 31580
rect 27672 31526 27674 31578
rect 27854 31526 27856 31578
rect 27610 31524 27616 31526
rect 27672 31524 27696 31526
rect 27752 31524 27776 31526
rect 27832 31524 27856 31526
rect 27912 31524 27918 31526
rect 27610 31515 27918 31524
rect 32610 31580 32918 31589
rect 32610 31578 32616 31580
rect 32672 31578 32696 31580
rect 32752 31578 32776 31580
rect 32832 31578 32856 31580
rect 32912 31578 32918 31580
rect 32672 31526 32674 31578
rect 32854 31526 32856 31578
rect 32610 31524 32616 31526
rect 32672 31524 32696 31526
rect 32752 31524 32776 31526
rect 32832 31524 32856 31526
rect 32912 31524 32918 31526
rect 32610 31515 32918 31524
rect 37610 31580 37918 31589
rect 37610 31578 37616 31580
rect 37672 31578 37696 31580
rect 37752 31578 37776 31580
rect 37832 31578 37856 31580
rect 37912 31578 37918 31580
rect 37672 31526 37674 31578
rect 37854 31526 37856 31578
rect 37610 31524 37616 31526
rect 37672 31524 37696 31526
rect 37752 31524 37776 31526
rect 37832 31524 37856 31526
rect 37912 31524 37918 31526
rect 37610 31515 37918 31524
rect 1950 31036 2258 31045
rect 1950 31034 1956 31036
rect 2012 31034 2036 31036
rect 2092 31034 2116 31036
rect 2172 31034 2196 31036
rect 2252 31034 2258 31036
rect 2012 30982 2014 31034
rect 2194 30982 2196 31034
rect 1950 30980 1956 30982
rect 2012 30980 2036 30982
rect 2092 30980 2116 30982
rect 2172 30980 2196 30982
rect 2252 30980 2258 30982
rect 1950 30971 2258 30980
rect 6950 31036 7258 31045
rect 6950 31034 6956 31036
rect 7012 31034 7036 31036
rect 7092 31034 7116 31036
rect 7172 31034 7196 31036
rect 7252 31034 7258 31036
rect 7012 30982 7014 31034
rect 7194 30982 7196 31034
rect 6950 30980 6956 30982
rect 7012 30980 7036 30982
rect 7092 30980 7116 30982
rect 7172 30980 7196 30982
rect 7252 30980 7258 30982
rect 6950 30971 7258 30980
rect 11950 31036 12258 31045
rect 11950 31034 11956 31036
rect 12012 31034 12036 31036
rect 12092 31034 12116 31036
rect 12172 31034 12196 31036
rect 12252 31034 12258 31036
rect 12012 30982 12014 31034
rect 12194 30982 12196 31034
rect 11950 30980 11956 30982
rect 12012 30980 12036 30982
rect 12092 30980 12116 30982
rect 12172 30980 12196 30982
rect 12252 30980 12258 30982
rect 11950 30971 12258 30980
rect 16950 31036 17258 31045
rect 16950 31034 16956 31036
rect 17012 31034 17036 31036
rect 17092 31034 17116 31036
rect 17172 31034 17196 31036
rect 17252 31034 17258 31036
rect 17012 30982 17014 31034
rect 17194 30982 17196 31034
rect 16950 30980 16956 30982
rect 17012 30980 17036 30982
rect 17092 30980 17116 30982
rect 17172 30980 17196 30982
rect 17252 30980 17258 30982
rect 16950 30971 17258 30980
rect 21950 31036 22258 31045
rect 21950 31034 21956 31036
rect 22012 31034 22036 31036
rect 22092 31034 22116 31036
rect 22172 31034 22196 31036
rect 22252 31034 22258 31036
rect 22012 30982 22014 31034
rect 22194 30982 22196 31034
rect 21950 30980 21956 30982
rect 22012 30980 22036 30982
rect 22092 30980 22116 30982
rect 22172 30980 22196 30982
rect 22252 30980 22258 30982
rect 21950 30971 22258 30980
rect 26950 31036 27258 31045
rect 26950 31034 26956 31036
rect 27012 31034 27036 31036
rect 27092 31034 27116 31036
rect 27172 31034 27196 31036
rect 27252 31034 27258 31036
rect 27012 30982 27014 31034
rect 27194 30982 27196 31034
rect 26950 30980 26956 30982
rect 27012 30980 27036 30982
rect 27092 30980 27116 30982
rect 27172 30980 27196 30982
rect 27252 30980 27258 30982
rect 26950 30971 27258 30980
rect 31950 31036 32258 31045
rect 31950 31034 31956 31036
rect 32012 31034 32036 31036
rect 32092 31034 32116 31036
rect 32172 31034 32196 31036
rect 32252 31034 32258 31036
rect 32012 30982 32014 31034
rect 32194 30982 32196 31034
rect 31950 30980 31956 30982
rect 32012 30980 32036 30982
rect 32092 30980 32116 30982
rect 32172 30980 32196 30982
rect 32252 30980 32258 30982
rect 31950 30971 32258 30980
rect 36950 31036 37258 31045
rect 36950 31034 36956 31036
rect 37012 31034 37036 31036
rect 37092 31034 37116 31036
rect 37172 31034 37196 31036
rect 37252 31034 37258 31036
rect 37012 30982 37014 31034
rect 37194 30982 37196 31034
rect 36950 30980 36956 30982
rect 37012 30980 37036 30982
rect 37092 30980 37116 30982
rect 37172 30980 37196 30982
rect 37252 30980 37258 30982
rect 36950 30971 37258 30980
rect 2610 30492 2918 30501
rect 2610 30490 2616 30492
rect 2672 30490 2696 30492
rect 2752 30490 2776 30492
rect 2832 30490 2856 30492
rect 2912 30490 2918 30492
rect 2672 30438 2674 30490
rect 2854 30438 2856 30490
rect 2610 30436 2616 30438
rect 2672 30436 2696 30438
rect 2752 30436 2776 30438
rect 2832 30436 2856 30438
rect 2912 30436 2918 30438
rect 2610 30427 2918 30436
rect 7610 30492 7918 30501
rect 7610 30490 7616 30492
rect 7672 30490 7696 30492
rect 7752 30490 7776 30492
rect 7832 30490 7856 30492
rect 7912 30490 7918 30492
rect 7672 30438 7674 30490
rect 7854 30438 7856 30490
rect 7610 30436 7616 30438
rect 7672 30436 7696 30438
rect 7752 30436 7776 30438
rect 7832 30436 7856 30438
rect 7912 30436 7918 30438
rect 7610 30427 7918 30436
rect 12610 30492 12918 30501
rect 12610 30490 12616 30492
rect 12672 30490 12696 30492
rect 12752 30490 12776 30492
rect 12832 30490 12856 30492
rect 12912 30490 12918 30492
rect 12672 30438 12674 30490
rect 12854 30438 12856 30490
rect 12610 30436 12616 30438
rect 12672 30436 12696 30438
rect 12752 30436 12776 30438
rect 12832 30436 12856 30438
rect 12912 30436 12918 30438
rect 12610 30427 12918 30436
rect 17610 30492 17918 30501
rect 17610 30490 17616 30492
rect 17672 30490 17696 30492
rect 17752 30490 17776 30492
rect 17832 30490 17856 30492
rect 17912 30490 17918 30492
rect 17672 30438 17674 30490
rect 17854 30438 17856 30490
rect 17610 30436 17616 30438
rect 17672 30436 17696 30438
rect 17752 30436 17776 30438
rect 17832 30436 17856 30438
rect 17912 30436 17918 30438
rect 17610 30427 17918 30436
rect 22610 30492 22918 30501
rect 22610 30490 22616 30492
rect 22672 30490 22696 30492
rect 22752 30490 22776 30492
rect 22832 30490 22856 30492
rect 22912 30490 22918 30492
rect 22672 30438 22674 30490
rect 22854 30438 22856 30490
rect 22610 30436 22616 30438
rect 22672 30436 22696 30438
rect 22752 30436 22776 30438
rect 22832 30436 22856 30438
rect 22912 30436 22918 30438
rect 22610 30427 22918 30436
rect 27610 30492 27918 30501
rect 27610 30490 27616 30492
rect 27672 30490 27696 30492
rect 27752 30490 27776 30492
rect 27832 30490 27856 30492
rect 27912 30490 27918 30492
rect 27672 30438 27674 30490
rect 27854 30438 27856 30490
rect 27610 30436 27616 30438
rect 27672 30436 27696 30438
rect 27752 30436 27776 30438
rect 27832 30436 27856 30438
rect 27912 30436 27918 30438
rect 27610 30427 27918 30436
rect 32610 30492 32918 30501
rect 32610 30490 32616 30492
rect 32672 30490 32696 30492
rect 32752 30490 32776 30492
rect 32832 30490 32856 30492
rect 32912 30490 32918 30492
rect 32672 30438 32674 30490
rect 32854 30438 32856 30490
rect 32610 30436 32616 30438
rect 32672 30436 32696 30438
rect 32752 30436 32776 30438
rect 32832 30436 32856 30438
rect 32912 30436 32918 30438
rect 32610 30427 32918 30436
rect 37610 30492 37918 30501
rect 37610 30490 37616 30492
rect 37672 30490 37696 30492
rect 37752 30490 37776 30492
rect 37832 30490 37856 30492
rect 37912 30490 37918 30492
rect 37672 30438 37674 30490
rect 37854 30438 37856 30490
rect 37610 30436 37616 30438
rect 37672 30436 37696 30438
rect 37752 30436 37776 30438
rect 37832 30436 37856 30438
rect 37912 30436 37918 30438
rect 37610 30427 37918 30436
rect 1950 29948 2258 29957
rect 1950 29946 1956 29948
rect 2012 29946 2036 29948
rect 2092 29946 2116 29948
rect 2172 29946 2196 29948
rect 2252 29946 2258 29948
rect 2012 29894 2014 29946
rect 2194 29894 2196 29946
rect 1950 29892 1956 29894
rect 2012 29892 2036 29894
rect 2092 29892 2116 29894
rect 2172 29892 2196 29894
rect 2252 29892 2258 29894
rect 1950 29883 2258 29892
rect 6950 29948 7258 29957
rect 6950 29946 6956 29948
rect 7012 29946 7036 29948
rect 7092 29946 7116 29948
rect 7172 29946 7196 29948
rect 7252 29946 7258 29948
rect 7012 29894 7014 29946
rect 7194 29894 7196 29946
rect 6950 29892 6956 29894
rect 7012 29892 7036 29894
rect 7092 29892 7116 29894
rect 7172 29892 7196 29894
rect 7252 29892 7258 29894
rect 6950 29883 7258 29892
rect 11950 29948 12258 29957
rect 11950 29946 11956 29948
rect 12012 29946 12036 29948
rect 12092 29946 12116 29948
rect 12172 29946 12196 29948
rect 12252 29946 12258 29948
rect 12012 29894 12014 29946
rect 12194 29894 12196 29946
rect 11950 29892 11956 29894
rect 12012 29892 12036 29894
rect 12092 29892 12116 29894
rect 12172 29892 12196 29894
rect 12252 29892 12258 29894
rect 11950 29883 12258 29892
rect 16950 29948 17258 29957
rect 16950 29946 16956 29948
rect 17012 29946 17036 29948
rect 17092 29946 17116 29948
rect 17172 29946 17196 29948
rect 17252 29946 17258 29948
rect 17012 29894 17014 29946
rect 17194 29894 17196 29946
rect 16950 29892 16956 29894
rect 17012 29892 17036 29894
rect 17092 29892 17116 29894
rect 17172 29892 17196 29894
rect 17252 29892 17258 29894
rect 16950 29883 17258 29892
rect 21950 29948 22258 29957
rect 21950 29946 21956 29948
rect 22012 29946 22036 29948
rect 22092 29946 22116 29948
rect 22172 29946 22196 29948
rect 22252 29946 22258 29948
rect 22012 29894 22014 29946
rect 22194 29894 22196 29946
rect 21950 29892 21956 29894
rect 22012 29892 22036 29894
rect 22092 29892 22116 29894
rect 22172 29892 22196 29894
rect 22252 29892 22258 29894
rect 21950 29883 22258 29892
rect 26950 29948 27258 29957
rect 26950 29946 26956 29948
rect 27012 29946 27036 29948
rect 27092 29946 27116 29948
rect 27172 29946 27196 29948
rect 27252 29946 27258 29948
rect 27012 29894 27014 29946
rect 27194 29894 27196 29946
rect 26950 29892 26956 29894
rect 27012 29892 27036 29894
rect 27092 29892 27116 29894
rect 27172 29892 27196 29894
rect 27252 29892 27258 29894
rect 26950 29883 27258 29892
rect 31950 29948 32258 29957
rect 31950 29946 31956 29948
rect 32012 29946 32036 29948
rect 32092 29946 32116 29948
rect 32172 29946 32196 29948
rect 32252 29946 32258 29948
rect 32012 29894 32014 29946
rect 32194 29894 32196 29946
rect 31950 29892 31956 29894
rect 32012 29892 32036 29894
rect 32092 29892 32116 29894
rect 32172 29892 32196 29894
rect 32252 29892 32258 29894
rect 31950 29883 32258 29892
rect 36950 29948 37258 29957
rect 36950 29946 36956 29948
rect 37012 29946 37036 29948
rect 37092 29946 37116 29948
rect 37172 29946 37196 29948
rect 37252 29946 37258 29948
rect 37012 29894 37014 29946
rect 37194 29894 37196 29946
rect 36950 29892 36956 29894
rect 37012 29892 37036 29894
rect 37092 29892 37116 29894
rect 37172 29892 37196 29894
rect 37252 29892 37258 29894
rect 36950 29883 37258 29892
rect 2610 29404 2918 29413
rect 2610 29402 2616 29404
rect 2672 29402 2696 29404
rect 2752 29402 2776 29404
rect 2832 29402 2856 29404
rect 2912 29402 2918 29404
rect 2672 29350 2674 29402
rect 2854 29350 2856 29402
rect 2610 29348 2616 29350
rect 2672 29348 2696 29350
rect 2752 29348 2776 29350
rect 2832 29348 2856 29350
rect 2912 29348 2918 29350
rect 2610 29339 2918 29348
rect 7610 29404 7918 29413
rect 7610 29402 7616 29404
rect 7672 29402 7696 29404
rect 7752 29402 7776 29404
rect 7832 29402 7856 29404
rect 7912 29402 7918 29404
rect 7672 29350 7674 29402
rect 7854 29350 7856 29402
rect 7610 29348 7616 29350
rect 7672 29348 7696 29350
rect 7752 29348 7776 29350
rect 7832 29348 7856 29350
rect 7912 29348 7918 29350
rect 7610 29339 7918 29348
rect 12610 29404 12918 29413
rect 12610 29402 12616 29404
rect 12672 29402 12696 29404
rect 12752 29402 12776 29404
rect 12832 29402 12856 29404
rect 12912 29402 12918 29404
rect 12672 29350 12674 29402
rect 12854 29350 12856 29402
rect 12610 29348 12616 29350
rect 12672 29348 12696 29350
rect 12752 29348 12776 29350
rect 12832 29348 12856 29350
rect 12912 29348 12918 29350
rect 12610 29339 12918 29348
rect 17610 29404 17918 29413
rect 17610 29402 17616 29404
rect 17672 29402 17696 29404
rect 17752 29402 17776 29404
rect 17832 29402 17856 29404
rect 17912 29402 17918 29404
rect 17672 29350 17674 29402
rect 17854 29350 17856 29402
rect 17610 29348 17616 29350
rect 17672 29348 17696 29350
rect 17752 29348 17776 29350
rect 17832 29348 17856 29350
rect 17912 29348 17918 29350
rect 17610 29339 17918 29348
rect 22610 29404 22918 29413
rect 22610 29402 22616 29404
rect 22672 29402 22696 29404
rect 22752 29402 22776 29404
rect 22832 29402 22856 29404
rect 22912 29402 22918 29404
rect 22672 29350 22674 29402
rect 22854 29350 22856 29402
rect 22610 29348 22616 29350
rect 22672 29348 22696 29350
rect 22752 29348 22776 29350
rect 22832 29348 22856 29350
rect 22912 29348 22918 29350
rect 22610 29339 22918 29348
rect 27610 29404 27918 29413
rect 27610 29402 27616 29404
rect 27672 29402 27696 29404
rect 27752 29402 27776 29404
rect 27832 29402 27856 29404
rect 27912 29402 27918 29404
rect 27672 29350 27674 29402
rect 27854 29350 27856 29402
rect 27610 29348 27616 29350
rect 27672 29348 27696 29350
rect 27752 29348 27776 29350
rect 27832 29348 27856 29350
rect 27912 29348 27918 29350
rect 27610 29339 27918 29348
rect 32610 29404 32918 29413
rect 32610 29402 32616 29404
rect 32672 29402 32696 29404
rect 32752 29402 32776 29404
rect 32832 29402 32856 29404
rect 32912 29402 32918 29404
rect 32672 29350 32674 29402
rect 32854 29350 32856 29402
rect 32610 29348 32616 29350
rect 32672 29348 32696 29350
rect 32752 29348 32776 29350
rect 32832 29348 32856 29350
rect 32912 29348 32918 29350
rect 32610 29339 32918 29348
rect 37610 29404 37918 29413
rect 37610 29402 37616 29404
rect 37672 29402 37696 29404
rect 37752 29402 37776 29404
rect 37832 29402 37856 29404
rect 37912 29402 37918 29404
rect 37672 29350 37674 29402
rect 37854 29350 37856 29402
rect 37610 29348 37616 29350
rect 37672 29348 37696 29350
rect 37752 29348 37776 29350
rect 37832 29348 37856 29350
rect 37912 29348 37918 29350
rect 37610 29339 37918 29348
rect 1950 28860 2258 28869
rect 1950 28858 1956 28860
rect 2012 28858 2036 28860
rect 2092 28858 2116 28860
rect 2172 28858 2196 28860
rect 2252 28858 2258 28860
rect 2012 28806 2014 28858
rect 2194 28806 2196 28858
rect 1950 28804 1956 28806
rect 2012 28804 2036 28806
rect 2092 28804 2116 28806
rect 2172 28804 2196 28806
rect 2252 28804 2258 28806
rect 1950 28795 2258 28804
rect 6950 28860 7258 28869
rect 6950 28858 6956 28860
rect 7012 28858 7036 28860
rect 7092 28858 7116 28860
rect 7172 28858 7196 28860
rect 7252 28858 7258 28860
rect 7012 28806 7014 28858
rect 7194 28806 7196 28858
rect 6950 28804 6956 28806
rect 7012 28804 7036 28806
rect 7092 28804 7116 28806
rect 7172 28804 7196 28806
rect 7252 28804 7258 28806
rect 6950 28795 7258 28804
rect 11950 28860 12258 28869
rect 11950 28858 11956 28860
rect 12012 28858 12036 28860
rect 12092 28858 12116 28860
rect 12172 28858 12196 28860
rect 12252 28858 12258 28860
rect 12012 28806 12014 28858
rect 12194 28806 12196 28858
rect 11950 28804 11956 28806
rect 12012 28804 12036 28806
rect 12092 28804 12116 28806
rect 12172 28804 12196 28806
rect 12252 28804 12258 28806
rect 11950 28795 12258 28804
rect 16950 28860 17258 28869
rect 16950 28858 16956 28860
rect 17012 28858 17036 28860
rect 17092 28858 17116 28860
rect 17172 28858 17196 28860
rect 17252 28858 17258 28860
rect 17012 28806 17014 28858
rect 17194 28806 17196 28858
rect 16950 28804 16956 28806
rect 17012 28804 17036 28806
rect 17092 28804 17116 28806
rect 17172 28804 17196 28806
rect 17252 28804 17258 28806
rect 16950 28795 17258 28804
rect 21950 28860 22258 28869
rect 21950 28858 21956 28860
rect 22012 28858 22036 28860
rect 22092 28858 22116 28860
rect 22172 28858 22196 28860
rect 22252 28858 22258 28860
rect 22012 28806 22014 28858
rect 22194 28806 22196 28858
rect 21950 28804 21956 28806
rect 22012 28804 22036 28806
rect 22092 28804 22116 28806
rect 22172 28804 22196 28806
rect 22252 28804 22258 28806
rect 21950 28795 22258 28804
rect 26950 28860 27258 28869
rect 26950 28858 26956 28860
rect 27012 28858 27036 28860
rect 27092 28858 27116 28860
rect 27172 28858 27196 28860
rect 27252 28858 27258 28860
rect 27012 28806 27014 28858
rect 27194 28806 27196 28858
rect 26950 28804 26956 28806
rect 27012 28804 27036 28806
rect 27092 28804 27116 28806
rect 27172 28804 27196 28806
rect 27252 28804 27258 28806
rect 26950 28795 27258 28804
rect 31950 28860 32258 28869
rect 31950 28858 31956 28860
rect 32012 28858 32036 28860
rect 32092 28858 32116 28860
rect 32172 28858 32196 28860
rect 32252 28858 32258 28860
rect 32012 28806 32014 28858
rect 32194 28806 32196 28858
rect 31950 28804 31956 28806
rect 32012 28804 32036 28806
rect 32092 28804 32116 28806
rect 32172 28804 32196 28806
rect 32252 28804 32258 28806
rect 31950 28795 32258 28804
rect 36950 28860 37258 28869
rect 36950 28858 36956 28860
rect 37012 28858 37036 28860
rect 37092 28858 37116 28860
rect 37172 28858 37196 28860
rect 37252 28858 37258 28860
rect 37012 28806 37014 28858
rect 37194 28806 37196 28858
rect 36950 28804 36956 28806
rect 37012 28804 37036 28806
rect 37092 28804 37116 28806
rect 37172 28804 37196 28806
rect 37252 28804 37258 28806
rect 36950 28795 37258 28804
rect 2610 28316 2918 28325
rect 2610 28314 2616 28316
rect 2672 28314 2696 28316
rect 2752 28314 2776 28316
rect 2832 28314 2856 28316
rect 2912 28314 2918 28316
rect 2672 28262 2674 28314
rect 2854 28262 2856 28314
rect 2610 28260 2616 28262
rect 2672 28260 2696 28262
rect 2752 28260 2776 28262
rect 2832 28260 2856 28262
rect 2912 28260 2918 28262
rect 2610 28251 2918 28260
rect 7610 28316 7918 28325
rect 7610 28314 7616 28316
rect 7672 28314 7696 28316
rect 7752 28314 7776 28316
rect 7832 28314 7856 28316
rect 7912 28314 7918 28316
rect 7672 28262 7674 28314
rect 7854 28262 7856 28314
rect 7610 28260 7616 28262
rect 7672 28260 7696 28262
rect 7752 28260 7776 28262
rect 7832 28260 7856 28262
rect 7912 28260 7918 28262
rect 7610 28251 7918 28260
rect 12610 28316 12918 28325
rect 12610 28314 12616 28316
rect 12672 28314 12696 28316
rect 12752 28314 12776 28316
rect 12832 28314 12856 28316
rect 12912 28314 12918 28316
rect 12672 28262 12674 28314
rect 12854 28262 12856 28314
rect 12610 28260 12616 28262
rect 12672 28260 12696 28262
rect 12752 28260 12776 28262
rect 12832 28260 12856 28262
rect 12912 28260 12918 28262
rect 12610 28251 12918 28260
rect 17610 28316 17918 28325
rect 17610 28314 17616 28316
rect 17672 28314 17696 28316
rect 17752 28314 17776 28316
rect 17832 28314 17856 28316
rect 17912 28314 17918 28316
rect 17672 28262 17674 28314
rect 17854 28262 17856 28314
rect 17610 28260 17616 28262
rect 17672 28260 17696 28262
rect 17752 28260 17776 28262
rect 17832 28260 17856 28262
rect 17912 28260 17918 28262
rect 17610 28251 17918 28260
rect 22610 28316 22918 28325
rect 22610 28314 22616 28316
rect 22672 28314 22696 28316
rect 22752 28314 22776 28316
rect 22832 28314 22856 28316
rect 22912 28314 22918 28316
rect 22672 28262 22674 28314
rect 22854 28262 22856 28314
rect 22610 28260 22616 28262
rect 22672 28260 22696 28262
rect 22752 28260 22776 28262
rect 22832 28260 22856 28262
rect 22912 28260 22918 28262
rect 22610 28251 22918 28260
rect 27610 28316 27918 28325
rect 27610 28314 27616 28316
rect 27672 28314 27696 28316
rect 27752 28314 27776 28316
rect 27832 28314 27856 28316
rect 27912 28314 27918 28316
rect 27672 28262 27674 28314
rect 27854 28262 27856 28314
rect 27610 28260 27616 28262
rect 27672 28260 27696 28262
rect 27752 28260 27776 28262
rect 27832 28260 27856 28262
rect 27912 28260 27918 28262
rect 27610 28251 27918 28260
rect 32610 28316 32918 28325
rect 32610 28314 32616 28316
rect 32672 28314 32696 28316
rect 32752 28314 32776 28316
rect 32832 28314 32856 28316
rect 32912 28314 32918 28316
rect 32672 28262 32674 28314
rect 32854 28262 32856 28314
rect 32610 28260 32616 28262
rect 32672 28260 32696 28262
rect 32752 28260 32776 28262
rect 32832 28260 32856 28262
rect 32912 28260 32918 28262
rect 32610 28251 32918 28260
rect 37610 28316 37918 28325
rect 37610 28314 37616 28316
rect 37672 28314 37696 28316
rect 37752 28314 37776 28316
rect 37832 28314 37856 28316
rect 37912 28314 37918 28316
rect 37672 28262 37674 28314
rect 37854 28262 37856 28314
rect 37610 28260 37616 28262
rect 37672 28260 37696 28262
rect 37752 28260 37776 28262
rect 37832 28260 37856 28262
rect 37912 28260 37918 28262
rect 37610 28251 37918 28260
rect 1950 27772 2258 27781
rect 1950 27770 1956 27772
rect 2012 27770 2036 27772
rect 2092 27770 2116 27772
rect 2172 27770 2196 27772
rect 2252 27770 2258 27772
rect 2012 27718 2014 27770
rect 2194 27718 2196 27770
rect 1950 27716 1956 27718
rect 2012 27716 2036 27718
rect 2092 27716 2116 27718
rect 2172 27716 2196 27718
rect 2252 27716 2258 27718
rect 1950 27707 2258 27716
rect 6950 27772 7258 27781
rect 6950 27770 6956 27772
rect 7012 27770 7036 27772
rect 7092 27770 7116 27772
rect 7172 27770 7196 27772
rect 7252 27770 7258 27772
rect 7012 27718 7014 27770
rect 7194 27718 7196 27770
rect 6950 27716 6956 27718
rect 7012 27716 7036 27718
rect 7092 27716 7116 27718
rect 7172 27716 7196 27718
rect 7252 27716 7258 27718
rect 6950 27707 7258 27716
rect 11950 27772 12258 27781
rect 11950 27770 11956 27772
rect 12012 27770 12036 27772
rect 12092 27770 12116 27772
rect 12172 27770 12196 27772
rect 12252 27770 12258 27772
rect 12012 27718 12014 27770
rect 12194 27718 12196 27770
rect 11950 27716 11956 27718
rect 12012 27716 12036 27718
rect 12092 27716 12116 27718
rect 12172 27716 12196 27718
rect 12252 27716 12258 27718
rect 11950 27707 12258 27716
rect 16950 27772 17258 27781
rect 16950 27770 16956 27772
rect 17012 27770 17036 27772
rect 17092 27770 17116 27772
rect 17172 27770 17196 27772
rect 17252 27770 17258 27772
rect 17012 27718 17014 27770
rect 17194 27718 17196 27770
rect 16950 27716 16956 27718
rect 17012 27716 17036 27718
rect 17092 27716 17116 27718
rect 17172 27716 17196 27718
rect 17252 27716 17258 27718
rect 16950 27707 17258 27716
rect 21950 27772 22258 27781
rect 21950 27770 21956 27772
rect 22012 27770 22036 27772
rect 22092 27770 22116 27772
rect 22172 27770 22196 27772
rect 22252 27770 22258 27772
rect 22012 27718 22014 27770
rect 22194 27718 22196 27770
rect 21950 27716 21956 27718
rect 22012 27716 22036 27718
rect 22092 27716 22116 27718
rect 22172 27716 22196 27718
rect 22252 27716 22258 27718
rect 21950 27707 22258 27716
rect 26950 27772 27258 27781
rect 26950 27770 26956 27772
rect 27012 27770 27036 27772
rect 27092 27770 27116 27772
rect 27172 27770 27196 27772
rect 27252 27770 27258 27772
rect 27012 27718 27014 27770
rect 27194 27718 27196 27770
rect 26950 27716 26956 27718
rect 27012 27716 27036 27718
rect 27092 27716 27116 27718
rect 27172 27716 27196 27718
rect 27252 27716 27258 27718
rect 26950 27707 27258 27716
rect 31950 27772 32258 27781
rect 31950 27770 31956 27772
rect 32012 27770 32036 27772
rect 32092 27770 32116 27772
rect 32172 27770 32196 27772
rect 32252 27770 32258 27772
rect 32012 27718 32014 27770
rect 32194 27718 32196 27770
rect 31950 27716 31956 27718
rect 32012 27716 32036 27718
rect 32092 27716 32116 27718
rect 32172 27716 32196 27718
rect 32252 27716 32258 27718
rect 31950 27707 32258 27716
rect 36950 27772 37258 27781
rect 36950 27770 36956 27772
rect 37012 27770 37036 27772
rect 37092 27770 37116 27772
rect 37172 27770 37196 27772
rect 37252 27770 37258 27772
rect 37012 27718 37014 27770
rect 37194 27718 37196 27770
rect 36950 27716 36956 27718
rect 37012 27716 37036 27718
rect 37092 27716 37116 27718
rect 37172 27716 37196 27718
rect 37252 27716 37258 27718
rect 36950 27707 37258 27716
rect 2610 27228 2918 27237
rect 2610 27226 2616 27228
rect 2672 27226 2696 27228
rect 2752 27226 2776 27228
rect 2832 27226 2856 27228
rect 2912 27226 2918 27228
rect 2672 27174 2674 27226
rect 2854 27174 2856 27226
rect 2610 27172 2616 27174
rect 2672 27172 2696 27174
rect 2752 27172 2776 27174
rect 2832 27172 2856 27174
rect 2912 27172 2918 27174
rect 2610 27163 2918 27172
rect 7610 27228 7918 27237
rect 7610 27226 7616 27228
rect 7672 27226 7696 27228
rect 7752 27226 7776 27228
rect 7832 27226 7856 27228
rect 7912 27226 7918 27228
rect 7672 27174 7674 27226
rect 7854 27174 7856 27226
rect 7610 27172 7616 27174
rect 7672 27172 7696 27174
rect 7752 27172 7776 27174
rect 7832 27172 7856 27174
rect 7912 27172 7918 27174
rect 7610 27163 7918 27172
rect 12610 27228 12918 27237
rect 12610 27226 12616 27228
rect 12672 27226 12696 27228
rect 12752 27226 12776 27228
rect 12832 27226 12856 27228
rect 12912 27226 12918 27228
rect 12672 27174 12674 27226
rect 12854 27174 12856 27226
rect 12610 27172 12616 27174
rect 12672 27172 12696 27174
rect 12752 27172 12776 27174
rect 12832 27172 12856 27174
rect 12912 27172 12918 27174
rect 12610 27163 12918 27172
rect 17610 27228 17918 27237
rect 17610 27226 17616 27228
rect 17672 27226 17696 27228
rect 17752 27226 17776 27228
rect 17832 27226 17856 27228
rect 17912 27226 17918 27228
rect 17672 27174 17674 27226
rect 17854 27174 17856 27226
rect 17610 27172 17616 27174
rect 17672 27172 17696 27174
rect 17752 27172 17776 27174
rect 17832 27172 17856 27174
rect 17912 27172 17918 27174
rect 17610 27163 17918 27172
rect 22610 27228 22918 27237
rect 22610 27226 22616 27228
rect 22672 27226 22696 27228
rect 22752 27226 22776 27228
rect 22832 27226 22856 27228
rect 22912 27226 22918 27228
rect 22672 27174 22674 27226
rect 22854 27174 22856 27226
rect 22610 27172 22616 27174
rect 22672 27172 22696 27174
rect 22752 27172 22776 27174
rect 22832 27172 22856 27174
rect 22912 27172 22918 27174
rect 22610 27163 22918 27172
rect 27610 27228 27918 27237
rect 27610 27226 27616 27228
rect 27672 27226 27696 27228
rect 27752 27226 27776 27228
rect 27832 27226 27856 27228
rect 27912 27226 27918 27228
rect 27672 27174 27674 27226
rect 27854 27174 27856 27226
rect 27610 27172 27616 27174
rect 27672 27172 27696 27174
rect 27752 27172 27776 27174
rect 27832 27172 27856 27174
rect 27912 27172 27918 27174
rect 27610 27163 27918 27172
rect 32610 27228 32918 27237
rect 32610 27226 32616 27228
rect 32672 27226 32696 27228
rect 32752 27226 32776 27228
rect 32832 27226 32856 27228
rect 32912 27226 32918 27228
rect 32672 27174 32674 27226
rect 32854 27174 32856 27226
rect 32610 27172 32616 27174
rect 32672 27172 32696 27174
rect 32752 27172 32776 27174
rect 32832 27172 32856 27174
rect 32912 27172 32918 27174
rect 32610 27163 32918 27172
rect 37610 27228 37918 27237
rect 37610 27226 37616 27228
rect 37672 27226 37696 27228
rect 37752 27226 37776 27228
rect 37832 27226 37856 27228
rect 37912 27226 37918 27228
rect 37672 27174 37674 27226
rect 37854 27174 37856 27226
rect 37610 27172 37616 27174
rect 37672 27172 37696 27174
rect 37752 27172 37776 27174
rect 37832 27172 37856 27174
rect 37912 27172 37918 27174
rect 37610 27163 37918 27172
rect 1950 26684 2258 26693
rect 1950 26682 1956 26684
rect 2012 26682 2036 26684
rect 2092 26682 2116 26684
rect 2172 26682 2196 26684
rect 2252 26682 2258 26684
rect 2012 26630 2014 26682
rect 2194 26630 2196 26682
rect 1950 26628 1956 26630
rect 2012 26628 2036 26630
rect 2092 26628 2116 26630
rect 2172 26628 2196 26630
rect 2252 26628 2258 26630
rect 1950 26619 2258 26628
rect 6950 26684 7258 26693
rect 6950 26682 6956 26684
rect 7012 26682 7036 26684
rect 7092 26682 7116 26684
rect 7172 26682 7196 26684
rect 7252 26682 7258 26684
rect 7012 26630 7014 26682
rect 7194 26630 7196 26682
rect 6950 26628 6956 26630
rect 7012 26628 7036 26630
rect 7092 26628 7116 26630
rect 7172 26628 7196 26630
rect 7252 26628 7258 26630
rect 6950 26619 7258 26628
rect 11950 26684 12258 26693
rect 11950 26682 11956 26684
rect 12012 26682 12036 26684
rect 12092 26682 12116 26684
rect 12172 26682 12196 26684
rect 12252 26682 12258 26684
rect 12012 26630 12014 26682
rect 12194 26630 12196 26682
rect 11950 26628 11956 26630
rect 12012 26628 12036 26630
rect 12092 26628 12116 26630
rect 12172 26628 12196 26630
rect 12252 26628 12258 26630
rect 11950 26619 12258 26628
rect 16950 26684 17258 26693
rect 16950 26682 16956 26684
rect 17012 26682 17036 26684
rect 17092 26682 17116 26684
rect 17172 26682 17196 26684
rect 17252 26682 17258 26684
rect 17012 26630 17014 26682
rect 17194 26630 17196 26682
rect 16950 26628 16956 26630
rect 17012 26628 17036 26630
rect 17092 26628 17116 26630
rect 17172 26628 17196 26630
rect 17252 26628 17258 26630
rect 16950 26619 17258 26628
rect 21950 26684 22258 26693
rect 21950 26682 21956 26684
rect 22012 26682 22036 26684
rect 22092 26682 22116 26684
rect 22172 26682 22196 26684
rect 22252 26682 22258 26684
rect 22012 26630 22014 26682
rect 22194 26630 22196 26682
rect 21950 26628 21956 26630
rect 22012 26628 22036 26630
rect 22092 26628 22116 26630
rect 22172 26628 22196 26630
rect 22252 26628 22258 26630
rect 21950 26619 22258 26628
rect 26950 26684 27258 26693
rect 26950 26682 26956 26684
rect 27012 26682 27036 26684
rect 27092 26682 27116 26684
rect 27172 26682 27196 26684
rect 27252 26682 27258 26684
rect 27012 26630 27014 26682
rect 27194 26630 27196 26682
rect 26950 26628 26956 26630
rect 27012 26628 27036 26630
rect 27092 26628 27116 26630
rect 27172 26628 27196 26630
rect 27252 26628 27258 26630
rect 26950 26619 27258 26628
rect 31950 26684 32258 26693
rect 31950 26682 31956 26684
rect 32012 26682 32036 26684
rect 32092 26682 32116 26684
rect 32172 26682 32196 26684
rect 32252 26682 32258 26684
rect 32012 26630 32014 26682
rect 32194 26630 32196 26682
rect 31950 26628 31956 26630
rect 32012 26628 32036 26630
rect 32092 26628 32116 26630
rect 32172 26628 32196 26630
rect 32252 26628 32258 26630
rect 31950 26619 32258 26628
rect 36950 26684 37258 26693
rect 36950 26682 36956 26684
rect 37012 26682 37036 26684
rect 37092 26682 37116 26684
rect 37172 26682 37196 26684
rect 37252 26682 37258 26684
rect 37012 26630 37014 26682
rect 37194 26630 37196 26682
rect 36950 26628 36956 26630
rect 37012 26628 37036 26630
rect 37092 26628 37116 26630
rect 37172 26628 37196 26630
rect 37252 26628 37258 26630
rect 36950 26619 37258 26628
rect 2610 26140 2918 26149
rect 2610 26138 2616 26140
rect 2672 26138 2696 26140
rect 2752 26138 2776 26140
rect 2832 26138 2856 26140
rect 2912 26138 2918 26140
rect 2672 26086 2674 26138
rect 2854 26086 2856 26138
rect 2610 26084 2616 26086
rect 2672 26084 2696 26086
rect 2752 26084 2776 26086
rect 2832 26084 2856 26086
rect 2912 26084 2918 26086
rect 2610 26075 2918 26084
rect 7610 26140 7918 26149
rect 7610 26138 7616 26140
rect 7672 26138 7696 26140
rect 7752 26138 7776 26140
rect 7832 26138 7856 26140
rect 7912 26138 7918 26140
rect 7672 26086 7674 26138
rect 7854 26086 7856 26138
rect 7610 26084 7616 26086
rect 7672 26084 7696 26086
rect 7752 26084 7776 26086
rect 7832 26084 7856 26086
rect 7912 26084 7918 26086
rect 7610 26075 7918 26084
rect 12610 26140 12918 26149
rect 12610 26138 12616 26140
rect 12672 26138 12696 26140
rect 12752 26138 12776 26140
rect 12832 26138 12856 26140
rect 12912 26138 12918 26140
rect 12672 26086 12674 26138
rect 12854 26086 12856 26138
rect 12610 26084 12616 26086
rect 12672 26084 12696 26086
rect 12752 26084 12776 26086
rect 12832 26084 12856 26086
rect 12912 26084 12918 26086
rect 12610 26075 12918 26084
rect 17610 26140 17918 26149
rect 17610 26138 17616 26140
rect 17672 26138 17696 26140
rect 17752 26138 17776 26140
rect 17832 26138 17856 26140
rect 17912 26138 17918 26140
rect 17672 26086 17674 26138
rect 17854 26086 17856 26138
rect 17610 26084 17616 26086
rect 17672 26084 17696 26086
rect 17752 26084 17776 26086
rect 17832 26084 17856 26086
rect 17912 26084 17918 26086
rect 17610 26075 17918 26084
rect 22610 26140 22918 26149
rect 22610 26138 22616 26140
rect 22672 26138 22696 26140
rect 22752 26138 22776 26140
rect 22832 26138 22856 26140
rect 22912 26138 22918 26140
rect 22672 26086 22674 26138
rect 22854 26086 22856 26138
rect 22610 26084 22616 26086
rect 22672 26084 22696 26086
rect 22752 26084 22776 26086
rect 22832 26084 22856 26086
rect 22912 26084 22918 26086
rect 22610 26075 22918 26084
rect 27610 26140 27918 26149
rect 27610 26138 27616 26140
rect 27672 26138 27696 26140
rect 27752 26138 27776 26140
rect 27832 26138 27856 26140
rect 27912 26138 27918 26140
rect 27672 26086 27674 26138
rect 27854 26086 27856 26138
rect 27610 26084 27616 26086
rect 27672 26084 27696 26086
rect 27752 26084 27776 26086
rect 27832 26084 27856 26086
rect 27912 26084 27918 26086
rect 27610 26075 27918 26084
rect 32610 26140 32918 26149
rect 32610 26138 32616 26140
rect 32672 26138 32696 26140
rect 32752 26138 32776 26140
rect 32832 26138 32856 26140
rect 32912 26138 32918 26140
rect 32672 26086 32674 26138
rect 32854 26086 32856 26138
rect 32610 26084 32616 26086
rect 32672 26084 32696 26086
rect 32752 26084 32776 26086
rect 32832 26084 32856 26086
rect 32912 26084 32918 26086
rect 32610 26075 32918 26084
rect 37610 26140 37918 26149
rect 37610 26138 37616 26140
rect 37672 26138 37696 26140
rect 37752 26138 37776 26140
rect 37832 26138 37856 26140
rect 37912 26138 37918 26140
rect 37672 26086 37674 26138
rect 37854 26086 37856 26138
rect 37610 26084 37616 26086
rect 37672 26084 37696 26086
rect 37752 26084 37776 26086
rect 37832 26084 37856 26086
rect 37912 26084 37918 26086
rect 37610 26075 37918 26084
rect 1950 25596 2258 25605
rect 1950 25594 1956 25596
rect 2012 25594 2036 25596
rect 2092 25594 2116 25596
rect 2172 25594 2196 25596
rect 2252 25594 2258 25596
rect 2012 25542 2014 25594
rect 2194 25542 2196 25594
rect 1950 25540 1956 25542
rect 2012 25540 2036 25542
rect 2092 25540 2116 25542
rect 2172 25540 2196 25542
rect 2252 25540 2258 25542
rect 1950 25531 2258 25540
rect 6950 25596 7258 25605
rect 6950 25594 6956 25596
rect 7012 25594 7036 25596
rect 7092 25594 7116 25596
rect 7172 25594 7196 25596
rect 7252 25594 7258 25596
rect 7012 25542 7014 25594
rect 7194 25542 7196 25594
rect 6950 25540 6956 25542
rect 7012 25540 7036 25542
rect 7092 25540 7116 25542
rect 7172 25540 7196 25542
rect 7252 25540 7258 25542
rect 6950 25531 7258 25540
rect 11950 25596 12258 25605
rect 11950 25594 11956 25596
rect 12012 25594 12036 25596
rect 12092 25594 12116 25596
rect 12172 25594 12196 25596
rect 12252 25594 12258 25596
rect 12012 25542 12014 25594
rect 12194 25542 12196 25594
rect 11950 25540 11956 25542
rect 12012 25540 12036 25542
rect 12092 25540 12116 25542
rect 12172 25540 12196 25542
rect 12252 25540 12258 25542
rect 11950 25531 12258 25540
rect 16950 25596 17258 25605
rect 16950 25594 16956 25596
rect 17012 25594 17036 25596
rect 17092 25594 17116 25596
rect 17172 25594 17196 25596
rect 17252 25594 17258 25596
rect 17012 25542 17014 25594
rect 17194 25542 17196 25594
rect 16950 25540 16956 25542
rect 17012 25540 17036 25542
rect 17092 25540 17116 25542
rect 17172 25540 17196 25542
rect 17252 25540 17258 25542
rect 16950 25531 17258 25540
rect 21950 25596 22258 25605
rect 21950 25594 21956 25596
rect 22012 25594 22036 25596
rect 22092 25594 22116 25596
rect 22172 25594 22196 25596
rect 22252 25594 22258 25596
rect 22012 25542 22014 25594
rect 22194 25542 22196 25594
rect 21950 25540 21956 25542
rect 22012 25540 22036 25542
rect 22092 25540 22116 25542
rect 22172 25540 22196 25542
rect 22252 25540 22258 25542
rect 21950 25531 22258 25540
rect 26950 25596 27258 25605
rect 26950 25594 26956 25596
rect 27012 25594 27036 25596
rect 27092 25594 27116 25596
rect 27172 25594 27196 25596
rect 27252 25594 27258 25596
rect 27012 25542 27014 25594
rect 27194 25542 27196 25594
rect 26950 25540 26956 25542
rect 27012 25540 27036 25542
rect 27092 25540 27116 25542
rect 27172 25540 27196 25542
rect 27252 25540 27258 25542
rect 26950 25531 27258 25540
rect 31950 25596 32258 25605
rect 31950 25594 31956 25596
rect 32012 25594 32036 25596
rect 32092 25594 32116 25596
rect 32172 25594 32196 25596
rect 32252 25594 32258 25596
rect 32012 25542 32014 25594
rect 32194 25542 32196 25594
rect 31950 25540 31956 25542
rect 32012 25540 32036 25542
rect 32092 25540 32116 25542
rect 32172 25540 32196 25542
rect 32252 25540 32258 25542
rect 31950 25531 32258 25540
rect 36950 25596 37258 25605
rect 36950 25594 36956 25596
rect 37012 25594 37036 25596
rect 37092 25594 37116 25596
rect 37172 25594 37196 25596
rect 37252 25594 37258 25596
rect 37012 25542 37014 25594
rect 37194 25542 37196 25594
rect 36950 25540 36956 25542
rect 37012 25540 37036 25542
rect 37092 25540 37116 25542
rect 37172 25540 37196 25542
rect 37252 25540 37258 25542
rect 36950 25531 37258 25540
rect 2610 25052 2918 25061
rect 2610 25050 2616 25052
rect 2672 25050 2696 25052
rect 2752 25050 2776 25052
rect 2832 25050 2856 25052
rect 2912 25050 2918 25052
rect 2672 24998 2674 25050
rect 2854 24998 2856 25050
rect 2610 24996 2616 24998
rect 2672 24996 2696 24998
rect 2752 24996 2776 24998
rect 2832 24996 2856 24998
rect 2912 24996 2918 24998
rect 2610 24987 2918 24996
rect 7610 25052 7918 25061
rect 7610 25050 7616 25052
rect 7672 25050 7696 25052
rect 7752 25050 7776 25052
rect 7832 25050 7856 25052
rect 7912 25050 7918 25052
rect 7672 24998 7674 25050
rect 7854 24998 7856 25050
rect 7610 24996 7616 24998
rect 7672 24996 7696 24998
rect 7752 24996 7776 24998
rect 7832 24996 7856 24998
rect 7912 24996 7918 24998
rect 7610 24987 7918 24996
rect 12610 25052 12918 25061
rect 12610 25050 12616 25052
rect 12672 25050 12696 25052
rect 12752 25050 12776 25052
rect 12832 25050 12856 25052
rect 12912 25050 12918 25052
rect 12672 24998 12674 25050
rect 12854 24998 12856 25050
rect 12610 24996 12616 24998
rect 12672 24996 12696 24998
rect 12752 24996 12776 24998
rect 12832 24996 12856 24998
rect 12912 24996 12918 24998
rect 12610 24987 12918 24996
rect 17610 25052 17918 25061
rect 17610 25050 17616 25052
rect 17672 25050 17696 25052
rect 17752 25050 17776 25052
rect 17832 25050 17856 25052
rect 17912 25050 17918 25052
rect 17672 24998 17674 25050
rect 17854 24998 17856 25050
rect 17610 24996 17616 24998
rect 17672 24996 17696 24998
rect 17752 24996 17776 24998
rect 17832 24996 17856 24998
rect 17912 24996 17918 24998
rect 17610 24987 17918 24996
rect 22610 25052 22918 25061
rect 22610 25050 22616 25052
rect 22672 25050 22696 25052
rect 22752 25050 22776 25052
rect 22832 25050 22856 25052
rect 22912 25050 22918 25052
rect 22672 24998 22674 25050
rect 22854 24998 22856 25050
rect 22610 24996 22616 24998
rect 22672 24996 22696 24998
rect 22752 24996 22776 24998
rect 22832 24996 22856 24998
rect 22912 24996 22918 24998
rect 22610 24987 22918 24996
rect 27610 25052 27918 25061
rect 27610 25050 27616 25052
rect 27672 25050 27696 25052
rect 27752 25050 27776 25052
rect 27832 25050 27856 25052
rect 27912 25050 27918 25052
rect 27672 24998 27674 25050
rect 27854 24998 27856 25050
rect 27610 24996 27616 24998
rect 27672 24996 27696 24998
rect 27752 24996 27776 24998
rect 27832 24996 27856 24998
rect 27912 24996 27918 24998
rect 27610 24987 27918 24996
rect 32610 25052 32918 25061
rect 32610 25050 32616 25052
rect 32672 25050 32696 25052
rect 32752 25050 32776 25052
rect 32832 25050 32856 25052
rect 32912 25050 32918 25052
rect 32672 24998 32674 25050
rect 32854 24998 32856 25050
rect 32610 24996 32616 24998
rect 32672 24996 32696 24998
rect 32752 24996 32776 24998
rect 32832 24996 32856 24998
rect 32912 24996 32918 24998
rect 32610 24987 32918 24996
rect 37610 25052 37918 25061
rect 37610 25050 37616 25052
rect 37672 25050 37696 25052
rect 37752 25050 37776 25052
rect 37832 25050 37856 25052
rect 37912 25050 37918 25052
rect 37672 24998 37674 25050
rect 37854 24998 37856 25050
rect 37610 24996 37616 24998
rect 37672 24996 37696 24998
rect 37752 24996 37776 24998
rect 37832 24996 37856 24998
rect 37912 24996 37918 24998
rect 37610 24987 37918 24996
rect 1950 24508 2258 24517
rect 1950 24506 1956 24508
rect 2012 24506 2036 24508
rect 2092 24506 2116 24508
rect 2172 24506 2196 24508
rect 2252 24506 2258 24508
rect 2012 24454 2014 24506
rect 2194 24454 2196 24506
rect 1950 24452 1956 24454
rect 2012 24452 2036 24454
rect 2092 24452 2116 24454
rect 2172 24452 2196 24454
rect 2252 24452 2258 24454
rect 1950 24443 2258 24452
rect 6950 24508 7258 24517
rect 6950 24506 6956 24508
rect 7012 24506 7036 24508
rect 7092 24506 7116 24508
rect 7172 24506 7196 24508
rect 7252 24506 7258 24508
rect 7012 24454 7014 24506
rect 7194 24454 7196 24506
rect 6950 24452 6956 24454
rect 7012 24452 7036 24454
rect 7092 24452 7116 24454
rect 7172 24452 7196 24454
rect 7252 24452 7258 24454
rect 6950 24443 7258 24452
rect 11950 24508 12258 24517
rect 11950 24506 11956 24508
rect 12012 24506 12036 24508
rect 12092 24506 12116 24508
rect 12172 24506 12196 24508
rect 12252 24506 12258 24508
rect 12012 24454 12014 24506
rect 12194 24454 12196 24506
rect 11950 24452 11956 24454
rect 12012 24452 12036 24454
rect 12092 24452 12116 24454
rect 12172 24452 12196 24454
rect 12252 24452 12258 24454
rect 11950 24443 12258 24452
rect 16950 24508 17258 24517
rect 16950 24506 16956 24508
rect 17012 24506 17036 24508
rect 17092 24506 17116 24508
rect 17172 24506 17196 24508
rect 17252 24506 17258 24508
rect 17012 24454 17014 24506
rect 17194 24454 17196 24506
rect 16950 24452 16956 24454
rect 17012 24452 17036 24454
rect 17092 24452 17116 24454
rect 17172 24452 17196 24454
rect 17252 24452 17258 24454
rect 16950 24443 17258 24452
rect 21950 24508 22258 24517
rect 21950 24506 21956 24508
rect 22012 24506 22036 24508
rect 22092 24506 22116 24508
rect 22172 24506 22196 24508
rect 22252 24506 22258 24508
rect 22012 24454 22014 24506
rect 22194 24454 22196 24506
rect 21950 24452 21956 24454
rect 22012 24452 22036 24454
rect 22092 24452 22116 24454
rect 22172 24452 22196 24454
rect 22252 24452 22258 24454
rect 21950 24443 22258 24452
rect 26950 24508 27258 24517
rect 26950 24506 26956 24508
rect 27012 24506 27036 24508
rect 27092 24506 27116 24508
rect 27172 24506 27196 24508
rect 27252 24506 27258 24508
rect 27012 24454 27014 24506
rect 27194 24454 27196 24506
rect 26950 24452 26956 24454
rect 27012 24452 27036 24454
rect 27092 24452 27116 24454
rect 27172 24452 27196 24454
rect 27252 24452 27258 24454
rect 26950 24443 27258 24452
rect 31950 24508 32258 24517
rect 31950 24506 31956 24508
rect 32012 24506 32036 24508
rect 32092 24506 32116 24508
rect 32172 24506 32196 24508
rect 32252 24506 32258 24508
rect 32012 24454 32014 24506
rect 32194 24454 32196 24506
rect 31950 24452 31956 24454
rect 32012 24452 32036 24454
rect 32092 24452 32116 24454
rect 32172 24452 32196 24454
rect 32252 24452 32258 24454
rect 31950 24443 32258 24452
rect 36950 24508 37258 24517
rect 36950 24506 36956 24508
rect 37012 24506 37036 24508
rect 37092 24506 37116 24508
rect 37172 24506 37196 24508
rect 37252 24506 37258 24508
rect 37012 24454 37014 24506
rect 37194 24454 37196 24506
rect 36950 24452 36956 24454
rect 37012 24452 37036 24454
rect 37092 24452 37116 24454
rect 37172 24452 37196 24454
rect 37252 24452 37258 24454
rect 36950 24443 37258 24452
rect 2610 23964 2918 23973
rect 2610 23962 2616 23964
rect 2672 23962 2696 23964
rect 2752 23962 2776 23964
rect 2832 23962 2856 23964
rect 2912 23962 2918 23964
rect 2672 23910 2674 23962
rect 2854 23910 2856 23962
rect 2610 23908 2616 23910
rect 2672 23908 2696 23910
rect 2752 23908 2776 23910
rect 2832 23908 2856 23910
rect 2912 23908 2918 23910
rect 2610 23899 2918 23908
rect 7610 23964 7918 23973
rect 7610 23962 7616 23964
rect 7672 23962 7696 23964
rect 7752 23962 7776 23964
rect 7832 23962 7856 23964
rect 7912 23962 7918 23964
rect 7672 23910 7674 23962
rect 7854 23910 7856 23962
rect 7610 23908 7616 23910
rect 7672 23908 7696 23910
rect 7752 23908 7776 23910
rect 7832 23908 7856 23910
rect 7912 23908 7918 23910
rect 7610 23899 7918 23908
rect 12610 23964 12918 23973
rect 12610 23962 12616 23964
rect 12672 23962 12696 23964
rect 12752 23962 12776 23964
rect 12832 23962 12856 23964
rect 12912 23962 12918 23964
rect 12672 23910 12674 23962
rect 12854 23910 12856 23962
rect 12610 23908 12616 23910
rect 12672 23908 12696 23910
rect 12752 23908 12776 23910
rect 12832 23908 12856 23910
rect 12912 23908 12918 23910
rect 12610 23899 12918 23908
rect 17610 23964 17918 23973
rect 17610 23962 17616 23964
rect 17672 23962 17696 23964
rect 17752 23962 17776 23964
rect 17832 23962 17856 23964
rect 17912 23962 17918 23964
rect 17672 23910 17674 23962
rect 17854 23910 17856 23962
rect 17610 23908 17616 23910
rect 17672 23908 17696 23910
rect 17752 23908 17776 23910
rect 17832 23908 17856 23910
rect 17912 23908 17918 23910
rect 17610 23899 17918 23908
rect 22610 23964 22918 23973
rect 22610 23962 22616 23964
rect 22672 23962 22696 23964
rect 22752 23962 22776 23964
rect 22832 23962 22856 23964
rect 22912 23962 22918 23964
rect 22672 23910 22674 23962
rect 22854 23910 22856 23962
rect 22610 23908 22616 23910
rect 22672 23908 22696 23910
rect 22752 23908 22776 23910
rect 22832 23908 22856 23910
rect 22912 23908 22918 23910
rect 22610 23899 22918 23908
rect 27610 23964 27918 23973
rect 27610 23962 27616 23964
rect 27672 23962 27696 23964
rect 27752 23962 27776 23964
rect 27832 23962 27856 23964
rect 27912 23962 27918 23964
rect 27672 23910 27674 23962
rect 27854 23910 27856 23962
rect 27610 23908 27616 23910
rect 27672 23908 27696 23910
rect 27752 23908 27776 23910
rect 27832 23908 27856 23910
rect 27912 23908 27918 23910
rect 27610 23899 27918 23908
rect 32610 23964 32918 23973
rect 32610 23962 32616 23964
rect 32672 23962 32696 23964
rect 32752 23962 32776 23964
rect 32832 23962 32856 23964
rect 32912 23962 32918 23964
rect 32672 23910 32674 23962
rect 32854 23910 32856 23962
rect 32610 23908 32616 23910
rect 32672 23908 32696 23910
rect 32752 23908 32776 23910
rect 32832 23908 32856 23910
rect 32912 23908 32918 23910
rect 32610 23899 32918 23908
rect 37610 23964 37918 23973
rect 37610 23962 37616 23964
rect 37672 23962 37696 23964
rect 37752 23962 37776 23964
rect 37832 23962 37856 23964
rect 37912 23962 37918 23964
rect 37672 23910 37674 23962
rect 37854 23910 37856 23962
rect 37610 23908 37616 23910
rect 37672 23908 37696 23910
rect 37752 23908 37776 23910
rect 37832 23908 37856 23910
rect 37912 23908 37918 23910
rect 37610 23899 37918 23908
rect 1950 23420 2258 23429
rect 1950 23418 1956 23420
rect 2012 23418 2036 23420
rect 2092 23418 2116 23420
rect 2172 23418 2196 23420
rect 2252 23418 2258 23420
rect 2012 23366 2014 23418
rect 2194 23366 2196 23418
rect 1950 23364 1956 23366
rect 2012 23364 2036 23366
rect 2092 23364 2116 23366
rect 2172 23364 2196 23366
rect 2252 23364 2258 23366
rect 1950 23355 2258 23364
rect 6950 23420 7258 23429
rect 6950 23418 6956 23420
rect 7012 23418 7036 23420
rect 7092 23418 7116 23420
rect 7172 23418 7196 23420
rect 7252 23418 7258 23420
rect 7012 23366 7014 23418
rect 7194 23366 7196 23418
rect 6950 23364 6956 23366
rect 7012 23364 7036 23366
rect 7092 23364 7116 23366
rect 7172 23364 7196 23366
rect 7252 23364 7258 23366
rect 6950 23355 7258 23364
rect 11950 23420 12258 23429
rect 11950 23418 11956 23420
rect 12012 23418 12036 23420
rect 12092 23418 12116 23420
rect 12172 23418 12196 23420
rect 12252 23418 12258 23420
rect 12012 23366 12014 23418
rect 12194 23366 12196 23418
rect 11950 23364 11956 23366
rect 12012 23364 12036 23366
rect 12092 23364 12116 23366
rect 12172 23364 12196 23366
rect 12252 23364 12258 23366
rect 11950 23355 12258 23364
rect 16950 23420 17258 23429
rect 16950 23418 16956 23420
rect 17012 23418 17036 23420
rect 17092 23418 17116 23420
rect 17172 23418 17196 23420
rect 17252 23418 17258 23420
rect 17012 23366 17014 23418
rect 17194 23366 17196 23418
rect 16950 23364 16956 23366
rect 17012 23364 17036 23366
rect 17092 23364 17116 23366
rect 17172 23364 17196 23366
rect 17252 23364 17258 23366
rect 16950 23355 17258 23364
rect 21950 23420 22258 23429
rect 21950 23418 21956 23420
rect 22012 23418 22036 23420
rect 22092 23418 22116 23420
rect 22172 23418 22196 23420
rect 22252 23418 22258 23420
rect 22012 23366 22014 23418
rect 22194 23366 22196 23418
rect 21950 23364 21956 23366
rect 22012 23364 22036 23366
rect 22092 23364 22116 23366
rect 22172 23364 22196 23366
rect 22252 23364 22258 23366
rect 21950 23355 22258 23364
rect 26950 23420 27258 23429
rect 26950 23418 26956 23420
rect 27012 23418 27036 23420
rect 27092 23418 27116 23420
rect 27172 23418 27196 23420
rect 27252 23418 27258 23420
rect 27012 23366 27014 23418
rect 27194 23366 27196 23418
rect 26950 23364 26956 23366
rect 27012 23364 27036 23366
rect 27092 23364 27116 23366
rect 27172 23364 27196 23366
rect 27252 23364 27258 23366
rect 26950 23355 27258 23364
rect 31950 23420 32258 23429
rect 31950 23418 31956 23420
rect 32012 23418 32036 23420
rect 32092 23418 32116 23420
rect 32172 23418 32196 23420
rect 32252 23418 32258 23420
rect 32012 23366 32014 23418
rect 32194 23366 32196 23418
rect 31950 23364 31956 23366
rect 32012 23364 32036 23366
rect 32092 23364 32116 23366
rect 32172 23364 32196 23366
rect 32252 23364 32258 23366
rect 31950 23355 32258 23364
rect 36950 23420 37258 23429
rect 36950 23418 36956 23420
rect 37012 23418 37036 23420
rect 37092 23418 37116 23420
rect 37172 23418 37196 23420
rect 37252 23418 37258 23420
rect 37012 23366 37014 23418
rect 37194 23366 37196 23418
rect 36950 23364 36956 23366
rect 37012 23364 37036 23366
rect 37092 23364 37116 23366
rect 37172 23364 37196 23366
rect 37252 23364 37258 23366
rect 36950 23355 37258 23364
rect 2610 22876 2918 22885
rect 2610 22874 2616 22876
rect 2672 22874 2696 22876
rect 2752 22874 2776 22876
rect 2832 22874 2856 22876
rect 2912 22874 2918 22876
rect 2672 22822 2674 22874
rect 2854 22822 2856 22874
rect 2610 22820 2616 22822
rect 2672 22820 2696 22822
rect 2752 22820 2776 22822
rect 2832 22820 2856 22822
rect 2912 22820 2918 22822
rect 2610 22811 2918 22820
rect 7610 22876 7918 22885
rect 7610 22874 7616 22876
rect 7672 22874 7696 22876
rect 7752 22874 7776 22876
rect 7832 22874 7856 22876
rect 7912 22874 7918 22876
rect 7672 22822 7674 22874
rect 7854 22822 7856 22874
rect 7610 22820 7616 22822
rect 7672 22820 7696 22822
rect 7752 22820 7776 22822
rect 7832 22820 7856 22822
rect 7912 22820 7918 22822
rect 7610 22811 7918 22820
rect 12610 22876 12918 22885
rect 12610 22874 12616 22876
rect 12672 22874 12696 22876
rect 12752 22874 12776 22876
rect 12832 22874 12856 22876
rect 12912 22874 12918 22876
rect 12672 22822 12674 22874
rect 12854 22822 12856 22874
rect 12610 22820 12616 22822
rect 12672 22820 12696 22822
rect 12752 22820 12776 22822
rect 12832 22820 12856 22822
rect 12912 22820 12918 22822
rect 12610 22811 12918 22820
rect 17610 22876 17918 22885
rect 17610 22874 17616 22876
rect 17672 22874 17696 22876
rect 17752 22874 17776 22876
rect 17832 22874 17856 22876
rect 17912 22874 17918 22876
rect 17672 22822 17674 22874
rect 17854 22822 17856 22874
rect 17610 22820 17616 22822
rect 17672 22820 17696 22822
rect 17752 22820 17776 22822
rect 17832 22820 17856 22822
rect 17912 22820 17918 22822
rect 17610 22811 17918 22820
rect 22610 22876 22918 22885
rect 22610 22874 22616 22876
rect 22672 22874 22696 22876
rect 22752 22874 22776 22876
rect 22832 22874 22856 22876
rect 22912 22874 22918 22876
rect 22672 22822 22674 22874
rect 22854 22822 22856 22874
rect 22610 22820 22616 22822
rect 22672 22820 22696 22822
rect 22752 22820 22776 22822
rect 22832 22820 22856 22822
rect 22912 22820 22918 22822
rect 22610 22811 22918 22820
rect 27610 22876 27918 22885
rect 27610 22874 27616 22876
rect 27672 22874 27696 22876
rect 27752 22874 27776 22876
rect 27832 22874 27856 22876
rect 27912 22874 27918 22876
rect 27672 22822 27674 22874
rect 27854 22822 27856 22874
rect 27610 22820 27616 22822
rect 27672 22820 27696 22822
rect 27752 22820 27776 22822
rect 27832 22820 27856 22822
rect 27912 22820 27918 22822
rect 27610 22811 27918 22820
rect 32610 22876 32918 22885
rect 32610 22874 32616 22876
rect 32672 22874 32696 22876
rect 32752 22874 32776 22876
rect 32832 22874 32856 22876
rect 32912 22874 32918 22876
rect 32672 22822 32674 22874
rect 32854 22822 32856 22874
rect 32610 22820 32616 22822
rect 32672 22820 32696 22822
rect 32752 22820 32776 22822
rect 32832 22820 32856 22822
rect 32912 22820 32918 22822
rect 32610 22811 32918 22820
rect 37610 22876 37918 22885
rect 37610 22874 37616 22876
rect 37672 22874 37696 22876
rect 37752 22874 37776 22876
rect 37832 22874 37856 22876
rect 37912 22874 37918 22876
rect 37672 22822 37674 22874
rect 37854 22822 37856 22874
rect 37610 22820 37616 22822
rect 37672 22820 37696 22822
rect 37752 22820 37776 22822
rect 37832 22820 37856 22822
rect 37912 22820 37918 22822
rect 37610 22811 37918 22820
rect 1950 22332 2258 22341
rect 1950 22330 1956 22332
rect 2012 22330 2036 22332
rect 2092 22330 2116 22332
rect 2172 22330 2196 22332
rect 2252 22330 2258 22332
rect 2012 22278 2014 22330
rect 2194 22278 2196 22330
rect 1950 22276 1956 22278
rect 2012 22276 2036 22278
rect 2092 22276 2116 22278
rect 2172 22276 2196 22278
rect 2252 22276 2258 22278
rect 1950 22267 2258 22276
rect 6950 22332 7258 22341
rect 6950 22330 6956 22332
rect 7012 22330 7036 22332
rect 7092 22330 7116 22332
rect 7172 22330 7196 22332
rect 7252 22330 7258 22332
rect 7012 22278 7014 22330
rect 7194 22278 7196 22330
rect 6950 22276 6956 22278
rect 7012 22276 7036 22278
rect 7092 22276 7116 22278
rect 7172 22276 7196 22278
rect 7252 22276 7258 22278
rect 6950 22267 7258 22276
rect 11950 22332 12258 22341
rect 11950 22330 11956 22332
rect 12012 22330 12036 22332
rect 12092 22330 12116 22332
rect 12172 22330 12196 22332
rect 12252 22330 12258 22332
rect 12012 22278 12014 22330
rect 12194 22278 12196 22330
rect 11950 22276 11956 22278
rect 12012 22276 12036 22278
rect 12092 22276 12116 22278
rect 12172 22276 12196 22278
rect 12252 22276 12258 22278
rect 11950 22267 12258 22276
rect 16950 22332 17258 22341
rect 16950 22330 16956 22332
rect 17012 22330 17036 22332
rect 17092 22330 17116 22332
rect 17172 22330 17196 22332
rect 17252 22330 17258 22332
rect 17012 22278 17014 22330
rect 17194 22278 17196 22330
rect 16950 22276 16956 22278
rect 17012 22276 17036 22278
rect 17092 22276 17116 22278
rect 17172 22276 17196 22278
rect 17252 22276 17258 22278
rect 16950 22267 17258 22276
rect 21950 22332 22258 22341
rect 21950 22330 21956 22332
rect 22012 22330 22036 22332
rect 22092 22330 22116 22332
rect 22172 22330 22196 22332
rect 22252 22330 22258 22332
rect 22012 22278 22014 22330
rect 22194 22278 22196 22330
rect 21950 22276 21956 22278
rect 22012 22276 22036 22278
rect 22092 22276 22116 22278
rect 22172 22276 22196 22278
rect 22252 22276 22258 22278
rect 21950 22267 22258 22276
rect 26950 22332 27258 22341
rect 26950 22330 26956 22332
rect 27012 22330 27036 22332
rect 27092 22330 27116 22332
rect 27172 22330 27196 22332
rect 27252 22330 27258 22332
rect 27012 22278 27014 22330
rect 27194 22278 27196 22330
rect 26950 22276 26956 22278
rect 27012 22276 27036 22278
rect 27092 22276 27116 22278
rect 27172 22276 27196 22278
rect 27252 22276 27258 22278
rect 26950 22267 27258 22276
rect 31950 22332 32258 22341
rect 31950 22330 31956 22332
rect 32012 22330 32036 22332
rect 32092 22330 32116 22332
rect 32172 22330 32196 22332
rect 32252 22330 32258 22332
rect 32012 22278 32014 22330
rect 32194 22278 32196 22330
rect 31950 22276 31956 22278
rect 32012 22276 32036 22278
rect 32092 22276 32116 22278
rect 32172 22276 32196 22278
rect 32252 22276 32258 22278
rect 31950 22267 32258 22276
rect 36950 22332 37258 22341
rect 36950 22330 36956 22332
rect 37012 22330 37036 22332
rect 37092 22330 37116 22332
rect 37172 22330 37196 22332
rect 37252 22330 37258 22332
rect 37012 22278 37014 22330
rect 37194 22278 37196 22330
rect 36950 22276 36956 22278
rect 37012 22276 37036 22278
rect 37092 22276 37116 22278
rect 37172 22276 37196 22278
rect 37252 22276 37258 22278
rect 36950 22267 37258 22276
rect 37280 22024 37332 22030
rect 37280 21966 37332 21972
rect 2610 21788 2918 21797
rect 2610 21786 2616 21788
rect 2672 21786 2696 21788
rect 2752 21786 2776 21788
rect 2832 21786 2856 21788
rect 2912 21786 2918 21788
rect 2672 21734 2674 21786
rect 2854 21734 2856 21786
rect 2610 21732 2616 21734
rect 2672 21732 2696 21734
rect 2752 21732 2776 21734
rect 2832 21732 2856 21734
rect 2912 21732 2918 21734
rect 2610 21723 2918 21732
rect 7610 21788 7918 21797
rect 7610 21786 7616 21788
rect 7672 21786 7696 21788
rect 7752 21786 7776 21788
rect 7832 21786 7856 21788
rect 7912 21786 7918 21788
rect 7672 21734 7674 21786
rect 7854 21734 7856 21786
rect 7610 21732 7616 21734
rect 7672 21732 7696 21734
rect 7752 21732 7776 21734
rect 7832 21732 7856 21734
rect 7912 21732 7918 21734
rect 7610 21723 7918 21732
rect 12610 21788 12918 21797
rect 12610 21786 12616 21788
rect 12672 21786 12696 21788
rect 12752 21786 12776 21788
rect 12832 21786 12856 21788
rect 12912 21786 12918 21788
rect 12672 21734 12674 21786
rect 12854 21734 12856 21786
rect 12610 21732 12616 21734
rect 12672 21732 12696 21734
rect 12752 21732 12776 21734
rect 12832 21732 12856 21734
rect 12912 21732 12918 21734
rect 12610 21723 12918 21732
rect 17610 21788 17918 21797
rect 17610 21786 17616 21788
rect 17672 21786 17696 21788
rect 17752 21786 17776 21788
rect 17832 21786 17856 21788
rect 17912 21786 17918 21788
rect 17672 21734 17674 21786
rect 17854 21734 17856 21786
rect 17610 21732 17616 21734
rect 17672 21732 17696 21734
rect 17752 21732 17776 21734
rect 17832 21732 17856 21734
rect 17912 21732 17918 21734
rect 17610 21723 17918 21732
rect 22610 21788 22918 21797
rect 22610 21786 22616 21788
rect 22672 21786 22696 21788
rect 22752 21786 22776 21788
rect 22832 21786 22856 21788
rect 22912 21786 22918 21788
rect 22672 21734 22674 21786
rect 22854 21734 22856 21786
rect 22610 21732 22616 21734
rect 22672 21732 22696 21734
rect 22752 21732 22776 21734
rect 22832 21732 22856 21734
rect 22912 21732 22918 21734
rect 22610 21723 22918 21732
rect 27610 21788 27918 21797
rect 27610 21786 27616 21788
rect 27672 21786 27696 21788
rect 27752 21786 27776 21788
rect 27832 21786 27856 21788
rect 27912 21786 27918 21788
rect 27672 21734 27674 21786
rect 27854 21734 27856 21786
rect 27610 21732 27616 21734
rect 27672 21732 27696 21734
rect 27752 21732 27776 21734
rect 27832 21732 27856 21734
rect 27912 21732 27918 21734
rect 27610 21723 27918 21732
rect 32610 21788 32918 21797
rect 32610 21786 32616 21788
rect 32672 21786 32696 21788
rect 32752 21786 32776 21788
rect 32832 21786 32856 21788
rect 32912 21786 32918 21788
rect 32672 21734 32674 21786
rect 32854 21734 32856 21786
rect 32610 21732 32616 21734
rect 32672 21732 32696 21734
rect 32752 21732 32776 21734
rect 32832 21732 32856 21734
rect 32912 21732 32918 21734
rect 32610 21723 32918 21732
rect 940 21548 992 21554
rect 940 21490 992 21496
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 952 21185 980 21490
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 938 21176 994 21185
rect 1596 21146 1624 21286
rect 1950 21244 2258 21253
rect 1950 21242 1956 21244
rect 2012 21242 2036 21244
rect 2092 21242 2116 21244
rect 2172 21242 2196 21244
rect 2252 21242 2258 21244
rect 2012 21190 2014 21242
rect 2194 21190 2196 21242
rect 1950 21188 1956 21190
rect 2012 21188 2036 21190
rect 2092 21188 2116 21190
rect 2172 21188 2196 21190
rect 2252 21188 2258 21190
rect 1950 21179 2258 21188
rect 6950 21244 7258 21253
rect 6950 21242 6956 21244
rect 7012 21242 7036 21244
rect 7092 21242 7116 21244
rect 7172 21242 7196 21244
rect 7252 21242 7258 21244
rect 7012 21190 7014 21242
rect 7194 21190 7196 21242
rect 6950 21188 6956 21190
rect 7012 21188 7036 21190
rect 7092 21188 7116 21190
rect 7172 21188 7196 21190
rect 7252 21188 7258 21190
rect 6950 21179 7258 21188
rect 11950 21244 12258 21253
rect 11950 21242 11956 21244
rect 12012 21242 12036 21244
rect 12092 21242 12116 21244
rect 12172 21242 12196 21244
rect 12252 21242 12258 21244
rect 12012 21190 12014 21242
rect 12194 21190 12196 21242
rect 11950 21188 11956 21190
rect 12012 21188 12036 21190
rect 12092 21188 12116 21190
rect 12172 21188 12196 21190
rect 12252 21188 12258 21190
rect 11950 21179 12258 21188
rect 16950 21244 17258 21253
rect 16950 21242 16956 21244
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17252 21242 17258 21244
rect 17012 21190 17014 21242
rect 17194 21190 17196 21242
rect 16950 21188 16956 21190
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 17252 21188 17258 21190
rect 16950 21179 17258 21188
rect 938 21111 994 21120
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 1400 20800 1452 20806
rect 1400 20742 1452 20748
rect 1412 20641 1440 20742
rect 2610 20700 2918 20709
rect 2610 20698 2616 20700
rect 2672 20698 2696 20700
rect 2752 20698 2776 20700
rect 2832 20698 2856 20700
rect 2912 20698 2918 20700
rect 2672 20646 2674 20698
rect 2854 20646 2856 20698
rect 2610 20644 2616 20646
rect 2672 20644 2696 20646
rect 2752 20644 2776 20646
rect 2832 20644 2856 20646
rect 2912 20644 2918 20646
rect 1398 20632 1454 20641
rect 2610 20635 2918 20644
rect 7610 20700 7918 20709
rect 7610 20698 7616 20700
rect 7672 20698 7696 20700
rect 7752 20698 7776 20700
rect 7832 20698 7856 20700
rect 7912 20698 7918 20700
rect 7672 20646 7674 20698
rect 7854 20646 7856 20698
rect 7610 20644 7616 20646
rect 7672 20644 7696 20646
rect 7752 20644 7776 20646
rect 7832 20644 7856 20646
rect 7912 20644 7918 20646
rect 7610 20635 7918 20644
rect 12610 20700 12918 20709
rect 12610 20698 12616 20700
rect 12672 20698 12696 20700
rect 12752 20698 12776 20700
rect 12832 20698 12856 20700
rect 12912 20698 12918 20700
rect 12672 20646 12674 20698
rect 12854 20646 12856 20698
rect 12610 20644 12616 20646
rect 12672 20644 12696 20646
rect 12752 20644 12776 20646
rect 12832 20644 12856 20646
rect 12912 20644 12918 20646
rect 12610 20635 12918 20644
rect 15212 20602 15240 20878
rect 1398 20567 1454 20576
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 1950 20156 2258 20165
rect 1950 20154 1956 20156
rect 2012 20154 2036 20156
rect 2092 20154 2116 20156
rect 2172 20154 2196 20156
rect 2252 20154 2258 20156
rect 2012 20102 2014 20154
rect 2194 20102 2196 20154
rect 1950 20100 1956 20102
rect 2012 20100 2036 20102
rect 2092 20100 2116 20102
rect 2172 20100 2196 20102
rect 2252 20100 2258 20102
rect 1950 20091 2258 20100
rect 6950 20156 7258 20165
rect 6950 20154 6956 20156
rect 7012 20154 7036 20156
rect 7092 20154 7116 20156
rect 7172 20154 7196 20156
rect 7252 20154 7258 20156
rect 7012 20102 7014 20154
rect 7194 20102 7196 20154
rect 6950 20100 6956 20102
rect 7012 20100 7036 20102
rect 7092 20100 7116 20102
rect 7172 20100 7196 20102
rect 7252 20100 7258 20102
rect 6950 20091 7258 20100
rect 11950 20156 12258 20165
rect 11950 20154 11956 20156
rect 12012 20154 12036 20156
rect 12092 20154 12116 20156
rect 12172 20154 12196 20156
rect 12252 20154 12258 20156
rect 12012 20102 12014 20154
rect 12194 20102 12196 20154
rect 11950 20100 11956 20102
rect 12012 20100 12036 20102
rect 12092 20100 12116 20102
rect 12172 20100 12196 20102
rect 12252 20100 12258 20102
rect 11950 20091 12258 20100
rect 15304 19854 15332 21082
rect 19812 21010 19840 21286
rect 19800 21004 19852 21010
rect 19800 20946 19852 20952
rect 19708 20868 19760 20874
rect 19708 20810 19760 20816
rect 17610 20700 17918 20709
rect 17610 20698 17616 20700
rect 17672 20698 17696 20700
rect 17752 20698 17776 20700
rect 17832 20698 17856 20700
rect 17912 20698 17918 20700
rect 17672 20646 17674 20698
rect 17854 20646 17856 20698
rect 17610 20644 17616 20646
rect 17672 20644 17696 20646
rect 17752 20644 17776 20646
rect 17832 20644 17856 20646
rect 17912 20644 17918 20646
rect 17610 20635 17918 20644
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 16950 20156 17258 20165
rect 16950 20154 16956 20156
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17252 20154 17258 20156
rect 17012 20102 17014 20154
rect 17194 20102 17196 20154
rect 16950 20100 16956 20102
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 17252 20100 17258 20102
rect 16950 20091 17258 20100
rect 940 19848 992 19854
rect 938 19816 940 19825
rect 15292 19848 15344 19854
rect 992 19816 994 19825
rect 15292 19790 15344 19796
rect 938 19751 994 19760
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 2610 19612 2918 19621
rect 2610 19610 2616 19612
rect 2672 19610 2696 19612
rect 2752 19610 2776 19612
rect 2832 19610 2856 19612
rect 2912 19610 2918 19612
rect 2672 19558 2674 19610
rect 2854 19558 2856 19610
rect 2610 19556 2616 19558
rect 2672 19556 2696 19558
rect 2752 19556 2776 19558
rect 2832 19556 2856 19558
rect 2912 19556 2918 19558
rect 2610 19547 2918 19556
rect 7610 19612 7918 19621
rect 7610 19610 7616 19612
rect 7672 19610 7696 19612
rect 7752 19610 7776 19612
rect 7832 19610 7856 19612
rect 7912 19610 7918 19612
rect 7672 19558 7674 19610
rect 7854 19558 7856 19610
rect 7610 19556 7616 19558
rect 7672 19556 7696 19558
rect 7752 19556 7776 19558
rect 7832 19556 7856 19558
rect 7912 19556 7918 19558
rect 7610 19547 7918 19556
rect 12610 19612 12918 19621
rect 12610 19610 12616 19612
rect 12672 19610 12696 19612
rect 12752 19610 12776 19612
rect 12832 19610 12856 19612
rect 12912 19610 12918 19612
rect 12672 19558 12674 19610
rect 12854 19558 12856 19610
rect 12610 19556 12616 19558
rect 12672 19556 12696 19558
rect 12752 19556 12776 19558
rect 12832 19556 12856 19558
rect 12912 19556 12918 19558
rect 12610 19547 12918 19556
rect 17610 19612 17918 19621
rect 17610 19610 17616 19612
rect 17672 19610 17696 19612
rect 17752 19610 17776 19612
rect 17832 19610 17856 19612
rect 17912 19610 17918 19612
rect 17672 19558 17674 19610
rect 17854 19558 17856 19610
rect 17610 19556 17616 19558
rect 17672 19556 17696 19558
rect 17752 19556 17776 19558
rect 17832 19556 17856 19558
rect 17912 19556 17918 19558
rect 17610 19547 17918 19556
rect 1400 19168 1452 19174
rect 1398 19136 1400 19145
rect 1452 19136 1454 19145
rect 1398 19071 1454 19080
rect 1950 19068 2258 19077
rect 1950 19066 1956 19068
rect 2012 19066 2036 19068
rect 2092 19066 2116 19068
rect 2172 19066 2196 19068
rect 2252 19066 2258 19068
rect 2012 19014 2014 19066
rect 2194 19014 2196 19066
rect 1950 19012 1956 19014
rect 2012 19012 2036 19014
rect 2092 19012 2116 19014
rect 2172 19012 2196 19014
rect 2252 19012 2258 19014
rect 1950 19003 2258 19012
rect 6950 19068 7258 19077
rect 6950 19066 6956 19068
rect 7012 19066 7036 19068
rect 7092 19066 7116 19068
rect 7172 19066 7196 19068
rect 7252 19066 7258 19068
rect 7012 19014 7014 19066
rect 7194 19014 7196 19066
rect 6950 19012 6956 19014
rect 7012 19012 7036 19014
rect 7092 19012 7116 19014
rect 7172 19012 7196 19014
rect 7252 19012 7258 19014
rect 6950 19003 7258 19012
rect 11950 19068 12258 19077
rect 11950 19066 11956 19068
rect 12012 19066 12036 19068
rect 12092 19066 12116 19068
rect 12172 19066 12196 19068
rect 12252 19066 12258 19068
rect 12012 19014 12014 19066
rect 12194 19014 12196 19066
rect 11950 19012 11956 19014
rect 12012 19012 12036 19014
rect 12092 19012 12116 19014
rect 12172 19012 12196 19014
rect 12252 19012 12258 19014
rect 11950 19003 12258 19012
rect 16950 19068 17258 19077
rect 16950 19066 16956 19068
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17252 19066 17258 19068
rect 17012 19014 17014 19066
rect 17194 19014 17196 19066
rect 16950 19012 16956 19014
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 17252 19012 17258 19014
rect 16950 19003 17258 19012
rect 18616 18902 18644 19654
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18984 19417 19012 19450
rect 18970 19408 19026 19417
rect 19352 19378 19380 20266
rect 18970 19343 19026 19352
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 19444 18834 19472 20402
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19536 19990 19564 20334
rect 19720 20262 19748 20810
rect 19812 20602 19840 20946
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19524 19984 19576 19990
rect 19524 19926 19576 19932
rect 19524 19780 19576 19786
rect 19524 19722 19576 19728
rect 19536 19174 19564 19722
rect 19720 19718 19748 20198
rect 19812 19922 19840 20538
rect 19904 19990 19932 20878
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 20180 20466 20208 20742
rect 20272 20602 20300 20810
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 19800 19916 19852 19922
rect 19800 19858 19852 19864
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19720 19378 19748 19654
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19536 18766 19564 19110
rect 940 18760 992 18766
rect 940 18702 992 18708
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 952 18465 980 18702
rect 2610 18524 2918 18533
rect 2610 18522 2616 18524
rect 2672 18522 2696 18524
rect 2752 18522 2776 18524
rect 2832 18522 2856 18524
rect 2912 18522 2918 18524
rect 2672 18470 2674 18522
rect 2854 18470 2856 18522
rect 2610 18468 2616 18470
rect 2672 18468 2696 18470
rect 2752 18468 2776 18470
rect 2832 18468 2856 18470
rect 2912 18468 2918 18470
rect 938 18456 994 18465
rect 2610 18459 2918 18468
rect 7610 18524 7918 18533
rect 7610 18522 7616 18524
rect 7672 18522 7696 18524
rect 7752 18522 7776 18524
rect 7832 18522 7856 18524
rect 7912 18522 7918 18524
rect 7672 18470 7674 18522
rect 7854 18470 7856 18522
rect 7610 18468 7616 18470
rect 7672 18468 7696 18470
rect 7752 18468 7776 18470
rect 7832 18468 7856 18470
rect 7912 18468 7918 18470
rect 7610 18459 7918 18468
rect 12610 18524 12918 18533
rect 12610 18522 12616 18524
rect 12672 18522 12696 18524
rect 12752 18522 12776 18524
rect 12832 18522 12856 18524
rect 12912 18522 12918 18524
rect 12672 18470 12674 18522
rect 12854 18470 12856 18522
rect 12610 18468 12616 18470
rect 12672 18468 12696 18470
rect 12752 18468 12776 18470
rect 12832 18468 12856 18470
rect 12912 18468 12918 18470
rect 12610 18459 12918 18468
rect 17610 18524 17918 18533
rect 17610 18522 17616 18524
rect 17672 18522 17696 18524
rect 17752 18522 17776 18524
rect 17832 18522 17856 18524
rect 17912 18522 17918 18524
rect 17672 18470 17674 18522
rect 17854 18470 17856 18522
rect 17610 18468 17616 18470
rect 17672 18468 17696 18470
rect 17752 18468 17776 18470
rect 17832 18468 17856 18470
rect 17912 18468 17918 18470
rect 17610 18459 17918 18468
rect 938 18391 994 18400
rect 19536 18358 19564 18702
rect 19720 18698 19748 19314
rect 19812 19242 19840 19858
rect 19904 19378 19932 19926
rect 20180 19378 20208 20402
rect 20456 19718 20484 21490
rect 21950 21244 22258 21253
rect 21950 21242 21956 21244
rect 22012 21242 22036 21244
rect 22092 21242 22116 21244
rect 22172 21242 22196 21244
rect 22252 21242 22258 21244
rect 22012 21190 22014 21242
rect 22194 21190 22196 21242
rect 21950 21188 21956 21190
rect 22012 21188 22036 21190
rect 22092 21188 22116 21190
rect 22172 21188 22196 21190
rect 22252 21188 22258 21190
rect 21950 21179 22258 21188
rect 26950 21244 27258 21253
rect 26950 21242 26956 21244
rect 27012 21242 27036 21244
rect 27092 21242 27116 21244
rect 27172 21242 27196 21244
rect 27252 21242 27258 21244
rect 27012 21190 27014 21242
rect 27194 21190 27196 21242
rect 26950 21188 26956 21190
rect 27012 21188 27036 21190
rect 27092 21188 27116 21190
rect 27172 21188 27196 21190
rect 27252 21188 27258 21190
rect 26950 21179 27258 21188
rect 31950 21244 32258 21253
rect 31950 21242 31956 21244
rect 32012 21242 32036 21244
rect 32092 21242 32116 21244
rect 32172 21242 32196 21244
rect 32252 21242 32258 21244
rect 32012 21190 32014 21242
rect 32194 21190 32196 21242
rect 31950 21188 31956 21190
rect 32012 21188 32036 21190
rect 32092 21188 32116 21190
rect 32172 21188 32196 21190
rect 32252 21188 32258 21190
rect 31950 21179 32258 21188
rect 36950 21244 37258 21253
rect 36950 21242 36956 21244
rect 37012 21242 37036 21244
rect 37092 21242 37116 21244
rect 37172 21242 37196 21244
rect 37252 21242 37258 21244
rect 37012 21190 37014 21242
rect 37194 21190 37196 21242
rect 36950 21188 36956 21190
rect 37012 21188 37036 21190
rect 37092 21188 37116 21190
rect 37172 21188 37196 21190
rect 37252 21188 37258 21190
rect 36950 21179 37258 21188
rect 34520 20936 34572 20942
rect 34520 20878 34572 20884
rect 22610 20700 22918 20709
rect 22610 20698 22616 20700
rect 22672 20698 22696 20700
rect 22752 20698 22776 20700
rect 22832 20698 22856 20700
rect 22912 20698 22918 20700
rect 22672 20646 22674 20698
rect 22854 20646 22856 20698
rect 22610 20644 22616 20646
rect 22672 20644 22696 20646
rect 22752 20644 22776 20646
rect 22832 20644 22856 20646
rect 22912 20644 22918 20646
rect 22610 20635 22918 20644
rect 27610 20700 27918 20709
rect 27610 20698 27616 20700
rect 27672 20698 27696 20700
rect 27752 20698 27776 20700
rect 27832 20698 27856 20700
rect 27912 20698 27918 20700
rect 27672 20646 27674 20698
rect 27854 20646 27856 20698
rect 27610 20644 27616 20646
rect 27672 20644 27696 20646
rect 27752 20644 27776 20646
rect 27832 20644 27856 20646
rect 27912 20644 27918 20646
rect 27610 20635 27918 20644
rect 32610 20700 32918 20709
rect 32610 20698 32616 20700
rect 32672 20698 32696 20700
rect 32752 20698 32776 20700
rect 32832 20698 32856 20700
rect 32912 20698 32918 20700
rect 32672 20646 32674 20698
rect 32854 20646 32856 20698
rect 32610 20644 32616 20646
rect 32672 20644 32696 20646
rect 32752 20644 32776 20646
rect 32832 20644 32856 20646
rect 32912 20644 32918 20646
rect 32610 20635 32918 20644
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 19800 19236 19852 19242
rect 19800 19178 19852 19184
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19720 18426 19748 18634
rect 19904 18630 19932 19314
rect 20180 19174 20208 19314
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20364 18698 20392 19110
rect 20456 18834 20484 19654
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20640 18630 20668 19178
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19904 18290 19932 18566
rect 20640 18290 20668 18566
rect 20732 18426 20760 20402
rect 21950 20156 22258 20165
rect 21950 20154 21956 20156
rect 22012 20154 22036 20156
rect 22092 20154 22116 20156
rect 22172 20154 22196 20156
rect 22252 20154 22258 20156
rect 22012 20102 22014 20154
rect 22194 20102 22196 20154
rect 21950 20100 21956 20102
rect 22012 20100 22036 20102
rect 22092 20100 22116 20102
rect 22172 20100 22196 20102
rect 22252 20100 22258 20102
rect 21950 20091 22258 20100
rect 26950 20156 27258 20165
rect 26950 20154 26956 20156
rect 27012 20154 27036 20156
rect 27092 20154 27116 20156
rect 27172 20154 27196 20156
rect 27252 20154 27258 20156
rect 27012 20102 27014 20154
rect 27194 20102 27196 20154
rect 26950 20100 26956 20102
rect 27012 20100 27036 20102
rect 27092 20100 27116 20102
rect 27172 20100 27196 20102
rect 27252 20100 27258 20102
rect 26950 20091 27258 20100
rect 31950 20156 32258 20165
rect 31950 20154 31956 20156
rect 32012 20154 32036 20156
rect 32092 20154 32116 20156
rect 32172 20154 32196 20156
rect 32252 20154 32258 20156
rect 32012 20102 32014 20154
rect 32194 20102 32196 20154
rect 31950 20100 31956 20102
rect 32012 20100 32036 20102
rect 32092 20100 32116 20102
rect 32172 20100 32196 20102
rect 32252 20100 32258 20102
rect 31950 20091 32258 20100
rect 34532 19990 34560 20878
rect 37292 20262 37320 21966
rect 38476 21888 38528 21894
rect 38474 21856 38476 21865
rect 38528 21856 38530 21865
rect 37610 21788 37918 21797
rect 38474 21791 38530 21800
rect 37610 21786 37616 21788
rect 37672 21786 37696 21788
rect 37752 21786 37776 21788
rect 37832 21786 37856 21788
rect 37912 21786 37918 21788
rect 37672 21734 37674 21786
rect 37854 21734 37856 21786
rect 37610 21732 37616 21734
rect 37672 21732 37696 21734
rect 37752 21732 37776 21734
rect 37832 21732 37856 21734
rect 37912 21732 37918 21734
rect 37610 21723 37918 21732
rect 38292 21548 38344 21554
rect 38292 21490 38344 21496
rect 37610 20700 37918 20709
rect 37610 20698 37616 20700
rect 37672 20698 37696 20700
rect 37752 20698 37776 20700
rect 37832 20698 37856 20700
rect 37912 20698 37918 20700
rect 37672 20646 37674 20698
rect 37854 20646 37856 20698
rect 37610 20644 37616 20646
rect 37672 20644 37696 20646
rect 37752 20644 37776 20646
rect 37832 20644 37856 20646
rect 37912 20644 37918 20646
rect 37610 20635 37918 20644
rect 38304 20330 38332 21490
rect 38476 21344 38528 21350
rect 38476 21286 38528 21292
rect 38488 21185 38516 21286
rect 38474 21176 38530 21185
rect 38474 21111 38530 21120
rect 39028 20732 39080 20738
rect 39028 20674 39080 20680
rect 39040 20505 39068 20674
rect 39026 20496 39082 20505
rect 39026 20431 39082 20440
rect 38292 20324 38344 20330
rect 38292 20266 38344 20272
rect 37280 20256 37332 20262
rect 37280 20198 37332 20204
rect 36950 20156 37258 20165
rect 36950 20154 36956 20156
rect 37012 20154 37036 20156
rect 37092 20154 37116 20156
rect 37172 20154 37196 20156
rect 37252 20154 37258 20156
rect 37012 20102 37014 20154
rect 37194 20102 37196 20154
rect 36950 20100 36956 20102
rect 37012 20100 37036 20102
rect 37092 20100 37116 20102
rect 37172 20100 37196 20102
rect 37252 20100 37258 20102
rect 36950 20091 37258 20100
rect 34520 19984 34572 19990
rect 34520 19926 34572 19932
rect 38844 19984 38896 19990
rect 38844 19926 38896 19932
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 26240 19848 26292 19854
rect 38856 19825 38884 19926
rect 26240 19790 26292 19796
rect 38842 19816 38898 19825
rect 21732 19780 21784 19786
rect 21732 19722 21784 19728
rect 21744 19514 21772 19722
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21100 18630 21128 19314
rect 21950 19068 22258 19077
rect 21950 19066 21956 19068
rect 22012 19066 22036 19068
rect 22092 19066 22116 19068
rect 22172 19066 22196 19068
rect 22252 19066 22258 19068
rect 22012 19014 22014 19066
rect 22194 19014 22196 19066
rect 21950 19012 21956 19014
rect 22012 19012 22036 19014
rect 22092 19012 22116 19014
rect 22172 19012 22196 19014
rect 22252 19012 22258 19014
rect 21950 19003 22258 19012
rect 22296 18970 22324 19790
rect 22610 19612 22918 19621
rect 22610 19610 22616 19612
rect 22672 19610 22696 19612
rect 22752 19610 22776 19612
rect 22832 19610 22856 19612
rect 22912 19610 22918 19612
rect 22672 19558 22674 19610
rect 22854 19558 22856 19610
rect 22610 19556 22616 19558
rect 22672 19556 22696 19558
rect 22752 19556 22776 19558
rect 22832 19556 22856 19558
rect 22912 19556 22918 19558
rect 22610 19547 22918 19556
rect 26252 19446 26280 19790
rect 38842 19751 38898 19760
rect 37280 19712 37332 19718
rect 37280 19654 37332 19660
rect 27610 19612 27918 19621
rect 27610 19610 27616 19612
rect 27672 19610 27696 19612
rect 27752 19610 27776 19612
rect 27832 19610 27856 19612
rect 27912 19610 27918 19612
rect 27672 19558 27674 19610
rect 27854 19558 27856 19610
rect 27610 19556 27616 19558
rect 27672 19556 27696 19558
rect 27752 19556 27776 19558
rect 27832 19556 27856 19558
rect 27912 19556 27918 19558
rect 27610 19547 27918 19556
rect 32610 19612 32918 19621
rect 32610 19610 32616 19612
rect 32672 19610 32696 19612
rect 32752 19610 32776 19612
rect 32832 19610 32856 19612
rect 32912 19610 32918 19612
rect 32672 19558 32674 19610
rect 32854 19558 32856 19610
rect 32610 19556 32616 19558
rect 32672 19556 32696 19558
rect 32752 19556 32776 19558
rect 32832 19556 32856 19558
rect 32912 19556 32918 19558
rect 32610 19547 32918 19556
rect 31760 19508 31812 19514
rect 31760 19450 31812 19456
rect 26240 19440 26292 19446
rect 26240 19382 26292 19388
rect 26950 19068 27258 19077
rect 26950 19066 26956 19068
rect 27012 19066 27036 19068
rect 27092 19066 27116 19068
rect 27172 19066 27196 19068
rect 27252 19066 27258 19068
rect 27012 19014 27014 19066
rect 27194 19014 27196 19066
rect 26950 19012 26956 19014
rect 27012 19012 27036 19014
rect 27092 19012 27116 19014
rect 27172 19012 27196 19014
rect 27252 19012 27258 19014
rect 26950 19003 27258 19012
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 21100 18358 21128 18566
rect 22610 18524 22918 18533
rect 22610 18522 22616 18524
rect 22672 18522 22696 18524
rect 22752 18522 22776 18524
rect 22832 18522 22856 18524
rect 22912 18522 22918 18524
rect 22672 18470 22674 18522
rect 22854 18470 22856 18522
rect 22610 18468 22616 18470
rect 22672 18468 22696 18470
rect 22752 18468 22776 18470
rect 22832 18468 22856 18470
rect 22912 18468 22918 18470
rect 22610 18459 22918 18468
rect 27610 18524 27918 18533
rect 27610 18522 27616 18524
rect 27672 18522 27696 18524
rect 27752 18522 27776 18524
rect 27832 18522 27856 18524
rect 27912 18522 27918 18524
rect 27672 18470 27674 18522
rect 27854 18470 27856 18522
rect 27610 18468 27616 18470
rect 27672 18468 27696 18470
rect 27752 18468 27776 18470
rect 27832 18468 27856 18470
rect 27912 18468 27918 18470
rect 27610 18459 27918 18468
rect 21088 18352 21140 18358
rect 21088 18294 21140 18300
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 1950 17980 2258 17989
rect 1950 17978 1956 17980
rect 2012 17978 2036 17980
rect 2092 17978 2116 17980
rect 2172 17978 2196 17980
rect 2252 17978 2258 17980
rect 2012 17926 2014 17978
rect 2194 17926 2196 17978
rect 1950 17924 1956 17926
rect 2012 17924 2036 17926
rect 2092 17924 2116 17926
rect 2172 17924 2196 17926
rect 2252 17924 2258 17926
rect 1950 17915 2258 17924
rect 6950 17980 7258 17989
rect 6950 17978 6956 17980
rect 7012 17978 7036 17980
rect 7092 17978 7116 17980
rect 7172 17978 7196 17980
rect 7252 17978 7258 17980
rect 7012 17926 7014 17978
rect 7194 17926 7196 17978
rect 6950 17924 6956 17926
rect 7012 17924 7036 17926
rect 7092 17924 7116 17926
rect 7172 17924 7196 17926
rect 7252 17924 7258 17926
rect 6950 17915 7258 17924
rect 11950 17980 12258 17989
rect 11950 17978 11956 17980
rect 12012 17978 12036 17980
rect 12092 17978 12116 17980
rect 12172 17978 12196 17980
rect 12252 17978 12258 17980
rect 12012 17926 12014 17978
rect 12194 17926 12196 17978
rect 11950 17924 11956 17926
rect 12012 17924 12036 17926
rect 12092 17924 12116 17926
rect 12172 17924 12196 17926
rect 12252 17924 12258 17926
rect 11950 17915 12258 17924
rect 16950 17980 17258 17989
rect 16950 17978 16956 17980
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17252 17978 17258 17980
rect 17012 17926 17014 17978
rect 17194 17926 17196 17978
rect 16950 17924 16956 17926
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 17252 17924 17258 17926
rect 16950 17915 17258 17924
rect 21950 17980 22258 17989
rect 21950 17978 21956 17980
rect 22012 17978 22036 17980
rect 22092 17978 22116 17980
rect 22172 17978 22196 17980
rect 22252 17978 22258 17980
rect 22012 17926 22014 17978
rect 22194 17926 22196 17978
rect 21950 17924 21956 17926
rect 22012 17924 22036 17926
rect 22092 17924 22116 17926
rect 22172 17924 22196 17926
rect 22252 17924 22258 17926
rect 21950 17915 22258 17924
rect 26950 17980 27258 17989
rect 26950 17978 26956 17980
rect 27012 17978 27036 17980
rect 27092 17978 27116 17980
rect 27172 17978 27196 17980
rect 27252 17978 27258 17980
rect 27012 17926 27014 17978
rect 27194 17926 27196 17978
rect 26950 17924 26956 17926
rect 27012 17924 27036 17926
rect 27092 17924 27116 17926
rect 27172 17924 27196 17926
rect 27252 17924 27258 17926
rect 26950 17915 27258 17924
rect 31772 17882 31800 19450
rect 31950 19068 32258 19077
rect 31950 19066 31956 19068
rect 32012 19066 32036 19068
rect 32092 19066 32116 19068
rect 32172 19066 32196 19068
rect 32252 19066 32258 19068
rect 32012 19014 32014 19066
rect 32194 19014 32196 19066
rect 31950 19012 31956 19014
rect 32012 19012 32036 19014
rect 32092 19012 32116 19014
rect 32172 19012 32196 19014
rect 32252 19012 32258 19014
rect 31950 19003 32258 19012
rect 36950 19068 37258 19077
rect 36950 19066 36956 19068
rect 37012 19066 37036 19068
rect 37092 19066 37116 19068
rect 37172 19066 37196 19068
rect 37252 19066 37258 19068
rect 37012 19014 37014 19066
rect 37194 19014 37196 19066
rect 36950 19012 36956 19014
rect 37012 19012 37036 19014
rect 37092 19012 37116 19014
rect 37172 19012 37196 19014
rect 37252 19012 37258 19014
rect 36950 19003 37258 19012
rect 37292 18766 37320 19654
rect 37610 19612 37918 19621
rect 37610 19610 37616 19612
rect 37672 19610 37696 19612
rect 37752 19610 37776 19612
rect 37832 19610 37856 19612
rect 37912 19610 37918 19612
rect 37672 19558 37674 19610
rect 37854 19558 37856 19610
rect 37610 19556 37616 19558
rect 37672 19556 37696 19558
rect 37752 19556 37776 19558
rect 37832 19556 37856 19558
rect 37912 19556 37918 19558
rect 37610 19547 37918 19556
rect 38290 19408 38346 19417
rect 38290 19343 38292 19352
rect 38344 19343 38346 19352
rect 38292 19314 38344 19320
rect 38476 19168 38528 19174
rect 38474 19136 38476 19145
rect 38528 19136 38530 19145
rect 38474 19071 38530 19080
rect 37280 18760 37332 18766
rect 37280 18702 37332 18708
rect 38476 18624 38528 18630
rect 38476 18566 38528 18572
rect 32610 18524 32918 18533
rect 32610 18522 32616 18524
rect 32672 18522 32696 18524
rect 32752 18522 32776 18524
rect 32832 18522 32856 18524
rect 32912 18522 32918 18524
rect 32672 18470 32674 18522
rect 32854 18470 32856 18522
rect 32610 18468 32616 18470
rect 32672 18468 32696 18470
rect 32752 18468 32776 18470
rect 32832 18468 32856 18470
rect 32912 18468 32918 18470
rect 32610 18459 32918 18468
rect 37610 18524 37918 18533
rect 37610 18522 37616 18524
rect 37672 18522 37696 18524
rect 37752 18522 37776 18524
rect 37832 18522 37856 18524
rect 37912 18522 37918 18524
rect 37672 18470 37674 18522
rect 37854 18470 37856 18522
rect 37610 18468 37616 18470
rect 37672 18468 37696 18470
rect 37752 18468 37776 18470
rect 37832 18468 37856 18470
rect 37912 18468 37918 18470
rect 37610 18459 37918 18468
rect 38488 18465 38516 18566
rect 38474 18456 38530 18465
rect 38474 18391 38530 18400
rect 31950 17980 32258 17989
rect 31950 17978 31956 17980
rect 32012 17978 32036 17980
rect 32092 17978 32116 17980
rect 32172 17978 32196 17980
rect 32252 17978 32258 17980
rect 32012 17926 32014 17978
rect 32194 17926 32196 17978
rect 31950 17924 31956 17926
rect 32012 17924 32036 17926
rect 32092 17924 32116 17926
rect 32172 17924 32196 17926
rect 32252 17924 32258 17926
rect 31950 17915 32258 17924
rect 36950 17980 37258 17989
rect 36950 17978 36956 17980
rect 37012 17978 37036 17980
rect 37092 17978 37116 17980
rect 37172 17978 37196 17980
rect 37252 17978 37258 17980
rect 37012 17926 37014 17978
rect 37194 17926 37196 17978
rect 36950 17924 36956 17926
rect 37012 17924 37036 17926
rect 37092 17924 37116 17926
rect 37172 17924 37196 17926
rect 37252 17924 37258 17926
rect 36950 17915 37258 17924
rect 31760 17876 31812 17882
rect 31760 17818 31812 17824
rect 34520 17876 34572 17882
rect 34520 17818 34572 17824
rect 34532 17785 34560 17818
rect 34518 17776 34574 17785
rect 34518 17711 34574 17720
rect 2610 17436 2918 17445
rect 2610 17434 2616 17436
rect 2672 17434 2696 17436
rect 2752 17434 2776 17436
rect 2832 17434 2856 17436
rect 2912 17434 2918 17436
rect 2672 17382 2674 17434
rect 2854 17382 2856 17434
rect 2610 17380 2616 17382
rect 2672 17380 2696 17382
rect 2752 17380 2776 17382
rect 2832 17380 2856 17382
rect 2912 17380 2918 17382
rect 2610 17371 2918 17380
rect 7610 17436 7918 17445
rect 7610 17434 7616 17436
rect 7672 17434 7696 17436
rect 7752 17434 7776 17436
rect 7832 17434 7856 17436
rect 7912 17434 7918 17436
rect 7672 17382 7674 17434
rect 7854 17382 7856 17434
rect 7610 17380 7616 17382
rect 7672 17380 7696 17382
rect 7752 17380 7776 17382
rect 7832 17380 7856 17382
rect 7912 17380 7918 17382
rect 7610 17371 7918 17380
rect 12610 17436 12918 17445
rect 12610 17434 12616 17436
rect 12672 17434 12696 17436
rect 12752 17434 12776 17436
rect 12832 17434 12856 17436
rect 12912 17434 12918 17436
rect 12672 17382 12674 17434
rect 12854 17382 12856 17434
rect 12610 17380 12616 17382
rect 12672 17380 12696 17382
rect 12752 17380 12776 17382
rect 12832 17380 12856 17382
rect 12912 17380 12918 17382
rect 12610 17371 12918 17380
rect 17610 17436 17918 17445
rect 17610 17434 17616 17436
rect 17672 17434 17696 17436
rect 17752 17434 17776 17436
rect 17832 17434 17856 17436
rect 17912 17434 17918 17436
rect 17672 17382 17674 17434
rect 17854 17382 17856 17434
rect 17610 17380 17616 17382
rect 17672 17380 17696 17382
rect 17752 17380 17776 17382
rect 17832 17380 17856 17382
rect 17912 17380 17918 17382
rect 17610 17371 17918 17380
rect 22610 17436 22918 17445
rect 22610 17434 22616 17436
rect 22672 17434 22696 17436
rect 22752 17434 22776 17436
rect 22832 17434 22856 17436
rect 22912 17434 22918 17436
rect 22672 17382 22674 17434
rect 22854 17382 22856 17434
rect 22610 17380 22616 17382
rect 22672 17380 22696 17382
rect 22752 17380 22776 17382
rect 22832 17380 22856 17382
rect 22912 17380 22918 17382
rect 22610 17371 22918 17380
rect 27610 17436 27918 17445
rect 27610 17434 27616 17436
rect 27672 17434 27696 17436
rect 27752 17434 27776 17436
rect 27832 17434 27856 17436
rect 27912 17434 27918 17436
rect 27672 17382 27674 17434
rect 27854 17382 27856 17434
rect 27610 17380 27616 17382
rect 27672 17380 27696 17382
rect 27752 17380 27776 17382
rect 27832 17380 27856 17382
rect 27912 17380 27918 17382
rect 27610 17371 27918 17380
rect 32610 17436 32918 17445
rect 32610 17434 32616 17436
rect 32672 17434 32696 17436
rect 32752 17434 32776 17436
rect 32832 17434 32856 17436
rect 32912 17434 32918 17436
rect 32672 17382 32674 17434
rect 32854 17382 32856 17434
rect 32610 17380 32616 17382
rect 32672 17380 32696 17382
rect 32752 17380 32776 17382
rect 32832 17380 32856 17382
rect 32912 17380 32918 17382
rect 32610 17371 32918 17380
rect 37610 17436 37918 17445
rect 37610 17434 37616 17436
rect 37672 17434 37696 17436
rect 37752 17434 37776 17436
rect 37832 17434 37856 17436
rect 37912 17434 37918 17436
rect 37672 17382 37674 17434
rect 37854 17382 37856 17434
rect 37610 17380 37616 17382
rect 37672 17380 37696 17382
rect 37752 17380 37776 17382
rect 37832 17380 37856 17382
rect 37912 17380 37918 17382
rect 37610 17371 37918 17380
rect 1950 16892 2258 16901
rect 1950 16890 1956 16892
rect 2012 16890 2036 16892
rect 2092 16890 2116 16892
rect 2172 16890 2196 16892
rect 2252 16890 2258 16892
rect 2012 16838 2014 16890
rect 2194 16838 2196 16890
rect 1950 16836 1956 16838
rect 2012 16836 2036 16838
rect 2092 16836 2116 16838
rect 2172 16836 2196 16838
rect 2252 16836 2258 16838
rect 1950 16827 2258 16836
rect 6950 16892 7258 16901
rect 6950 16890 6956 16892
rect 7012 16890 7036 16892
rect 7092 16890 7116 16892
rect 7172 16890 7196 16892
rect 7252 16890 7258 16892
rect 7012 16838 7014 16890
rect 7194 16838 7196 16890
rect 6950 16836 6956 16838
rect 7012 16836 7036 16838
rect 7092 16836 7116 16838
rect 7172 16836 7196 16838
rect 7252 16836 7258 16838
rect 6950 16827 7258 16836
rect 11950 16892 12258 16901
rect 11950 16890 11956 16892
rect 12012 16890 12036 16892
rect 12092 16890 12116 16892
rect 12172 16890 12196 16892
rect 12252 16890 12258 16892
rect 12012 16838 12014 16890
rect 12194 16838 12196 16890
rect 11950 16836 11956 16838
rect 12012 16836 12036 16838
rect 12092 16836 12116 16838
rect 12172 16836 12196 16838
rect 12252 16836 12258 16838
rect 11950 16827 12258 16836
rect 16950 16892 17258 16901
rect 16950 16890 16956 16892
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17252 16890 17258 16892
rect 17012 16838 17014 16890
rect 17194 16838 17196 16890
rect 16950 16836 16956 16838
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 17252 16836 17258 16838
rect 16950 16827 17258 16836
rect 21950 16892 22258 16901
rect 21950 16890 21956 16892
rect 22012 16890 22036 16892
rect 22092 16890 22116 16892
rect 22172 16890 22196 16892
rect 22252 16890 22258 16892
rect 22012 16838 22014 16890
rect 22194 16838 22196 16890
rect 21950 16836 21956 16838
rect 22012 16836 22036 16838
rect 22092 16836 22116 16838
rect 22172 16836 22196 16838
rect 22252 16836 22258 16838
rect 21950 16827 22258 16836
rect 26950 16892 27258 16901
rect 26950 16890 26956 16892
rect 27012 16890 27036 16892
rect 27092 16890 27116 16892
rect 27172 16890 27196 16892
rect 27252 16890 27258 16892
rect 27012 16838 27014 16890
rect 27194 16838 27196 16890
rect 26950 16836 26956 16838
rect 27012 16836 27036 16838
rect 27092 16836 27116 16838
rect 27172 16836 27196 16838
rect 27252 16836 27258 16838
rect 26950 16827 27258 16836
rect 31950 16892 32258 16901
rect 31950 16890 31956 16892
rect 32012 16890 32036 16892
rect 32092 16890 32116 16892
rect 32172 16890 32196 16892
rect 32252 16890 32258 16892
rect 32012 16838 32014 16890
rect 32194 16838 32196 16890
rect 31950 16836 31956 16838
rect 32012 16836 32036 16838
rect 32092 16836 32116 16838
rect 32172 16836 32196 16838
rect 32252 16836 32258 16838
rect 31950 16827 32258 16836
rect 36950 16892 37258 16901
rect 36950 16890 36956 16892
rect 37012 16890 37036 16892
rect 37092 16890 37116 16892
rect 37172 16890 37196 16892
rect 37252 16890 37258 16892
rect 37012 16838 37014 16890
rect 37194 16838 37196 16890
rect 36950 16836 36956 16838
rect 37012 16836 37036 16838
rect 37092 16836 37116 16838
rect 37172 16836 37196 16838
rect 37252 16836 37258 16838
rect 36950 16827 37258 16836
rect 2610 16348 2918 16357
rect 2610 16346 2616 16348
rect 2672 16346 2696 16348
rect 2752 16346 2776 16348
rect 2832 16346 2856 16348
rect 2912 16346 2918 16348
rect 2672 16294 2674 16346
rect 2854 16294 2856 16346
rect 2610 16292 2616 16294
rect 2672 16292 2696 16294
rect 2752 16292 2776 16294
rect 2832 16292 2856 16294
rect 2912 16292 2918 16294
rect 2610 16283 2918 16292
rect 7610 16348 7918 16357
rect 7610 16346 7616 16348
rect 7672 16346 7696 16348
rect 7752 16346 7776 16348
rect 7832 16346 7856 16348
rect 7912 16346 7918 16348
rect 7672 16294 7674 16346
rect 7854 16294 7856 16346
rect 7610 16292 7616 16294
rect 7672 16292 7696 16294
rect 7752 16292 7776 16294
rect 7832 16292 7856 16294
rect 7912 16292 7918 16294
rect 7610 16283 7918 16292
rect 12610 16348 12918 16357
rect 12610 16346 12616 16348
rect 12672 16346 12696 16348
rect 12752 16346 12776 16348
rect 12832 16346 12856 16348
rect 12912 16346 12918 16348
rect 12672 16294 12674 16346
rect 12854 16294 12856 16346
rect 12610 16292 12616 16294
rect 12672 16292 12696 16294
rect 12752 16292 12776 16294
rect 12832 16292 12856 16294
rect 12912 16292 12918 16294
rect 12610 16283 12918 16292
rect 17610 16348 17918 16357
rect 17610 16346 17616 16348
rect 17672 16346 17696 16348
rect 17752 16346 17776 16348
rect 17832 16346 17856 16348
rect 17912 16346 17918 16348
rect 17672 16294 17674 16346
rect 17854 16294 17856 16346
rect 17610 16292 17616 16294
rect 17672 16292 17696 16294
rect 17752 16292 17776 16294
rect 17832 16292 17856 16294
rect 17912 16292 17918 16294
rect 17610 16283 17918 16292
rect 22610 16348 22918 16357
rect 22610 16346 22616 16348
rect 22672 16346 22696 16348
rect 22752 16346 22776 16348
rect 22832 16346 22856 16348
rect 22912 16346 22918 16348
rect 22672 16294 22674 16346
rect 22854 16294 22856 16346
rect 22610 16292 22616 16294
rect 22672 16292 22696 16294
rect 22752 16292 22776 16294
rect 22832 16292 22856 16294
rect 22912 16292 22918 16294
rect 22610 16283 22918 16292
rect 27610 16348 27918 16357
rect 27610 16346 27616 16348
rect 27672 16346 27696 16348
rect 27752 16346 27776 16348
rect 27832 16346 27856 16348
rect 27912 16346 27918 16348
rect 27672 16294 27674 16346
rect 27854 16294 27856 16346
rect 27610 16292 27616 16294
rect 27672 16292 27696 16294
rect 27752 16292 27776 16294
rect 27832 16292 27856 16294
rect 27912 16292 27918 16294
rect 27610 16283 27918 16292
rect 32610 16348 32918 16357
rect 32610 16346 32616 16348
rect 32672 16346 32696 16348
rect 32752 16346 32776 16348
rect 32832 16346 32856 16348
rect 32912 16346 32918 16348
rect 32672 16294 32674 16346
rect 32854 16294 32856 16346
rect 32610 16292 32616 16294
rect 32672 16292 32696 16294
rect 32752 16292 32776 16294
rect 32832 16292 32856 16294
rect 32912 16292 32918 16294
rect 32610 16283 32918 16292
rect 37610 16348 37918 16357
rect 37610 16346 37616 16348
rect 37672 16346 37696 16348
rect 37752 16346 37776 16348
rect 37832 16346 37856 16348
rect 37912 16346 37918 16348
rect 37672 16294 37674 16346
rect 37854 16294 37856 16346
rect 37610 16292 37616 16294
rect 37672 16292 37696 16294
rect 37752 16292 37776 16294
rect 37832 16292 37856 16294
rect 37912 16292 37918 16294
rect 37610 16283 37918 16292
rect 1950 15804 2258 15813
rect 1950 15802 1956 15804
rect 2012 15802 2036 15804
rect 2092 15802 2116 15804
rect 2172 15802 2196 15804
rect 2252 15802 2258 15804
rect 2012 15750 2014 15802
rect 2194 15750 2196 15802
rect 1950 15748 1956 15750
rect 2012 15748 2036 15750
rect 2092 15748 2116 15750
rect 2172 15748 2196 15750
rect 2252 15748 2258 15750
rect 1950 15739 2258 15748
rect 6950 15804 7258 15813
rect 6950 15802 6956 15804
rect 7012 15802 7036 15804
rect 7092 15802 7116 15804
rect 7172 15802 7196 15804
rect 7252 15802 7258 15804
rect 7012 15750 7014 15802
rect 7194 15750 7196 15802
rect 6950 15748 6956 15750
rect 7012 15748 7036 15750
rect 7092 15748 7116 15750
rect 7172 15748 7196 15750
rect 7252 15748 7258 15750
rect 6950 15739 7258 15748
rect 11950 15804 12258 15813
rect 11950 15802 11956 15804
rect 12012 15802 12036 15804
rect 12092 15802 12116 15804
rect 12172 15802 12196 15804
rect 12252 15802 12258 15804
rect 12012 15750 12014 15802
rect 12194 15750 12196 15802
rect 11950 15748 11956 15750
rect 12012 15748 12036 15750
rect 12092 15748 12116 15750
rect 12172 15748 12196 15750
rect 12252 15748 12258 15750
rect 11950 15739 12258 15748
rect 16950 15804 17258 15813
rect 16950 15802 16956 15804
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17252 15802 17258 15804
rect 17012 15750 17014 15802
rect 17194 15750 17196 15802
rect 16950 15748 16956 15750
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 17252 15748 17258 15750
rect 16950 15739 17258 15748
rect 21950 15804 22258 15813
rect 21950 15802 21956 15804
rect 22012 15802 22036 15804
rect 22092 15802 22116 15804
rect 22172 15802 22196 15804
rect 22252 15802 22258 15804
rect 22012 15750 22014 15802
rect 22194 15750 22196 15802
rect 21950 15748 21956 15750
rect 22012 15748 22036 15750
rect 22092 15748 22116 15750
rect 22172 15748 22196 15750
rect 22252 15748 22258 15750
rect 21950 15739 22258 15748
rect 26950 15804 27258 15813
rect 26950 15802 26956 15804
rect 27012 15802 27036 15804
rect 27092 15802 27116 15804
rect 27172 15802 27196 15804
rect 27252 15802 27258 15804
rect 27012 15750 27014 15802
rect 27194 15750 27196 15802
rect 26950 15748 26956 15750
rect 27012 15748 27036 15750
rect 27092 15748 27116 15750
rect 27172 15748 27196 15750
rect 27252 15748 27258 15750
rect 26950 15739 27258 15748
rect 31950 15804 32258 15813
rect 31950 15802 31956 15804
rect 32012 15802 32036 15804
rect 32092 15802 32116 15804
rect 32172 15802 32196 15804
rect 32252 15802 32258 15804
rect 32012 15750 32014 15802
rect 32194 15750 32196 15802
rect 31950 15748 31956 15750
rect 32012 15748 32036 15750
rect 32092 15748 32116 15750
rect 32172 15748 32196 15750
rect 32252 15748 32258 15750
rect 31950 15739 32258 15748
rect 36950 15804 37258 15813
rect 36950 15802 36956 15804
rect 37012 15802 37036 15804
rect 37092 15802 37116 15804
rect 37172 15802 37196 15804
rect 37252 15802 37258 15804
rect 37012 15750 37014 15802
rect 37194 15750 37196 15802
rect 36950 15748 36956 15750
rect 37012 15748 37036 15750
rect 37092 15748 37116 15750
rect 37172 15748 37196 15750
rect 37252 15748 37258 15750
rect 36950 15739 37258 15748
rect 2610 15260 2918 15269
rect 2610 15258 2616 15260
rect 2672 15258 2696 15260
rect 2752 15258 2776 15260
rect 2832 15258 2856 15260
rect 2912 15258 2918 15260
rect 2672 15206 2674 15258
rect 2854 15206 2856 15258
rect 2610 15204 2616 15206
rect 2672 15204 2696 15206
rect 2752 15204 2776 15206
rect 2832 15204 2856 15206
rect 2912 15204 2918 15206
rect 2610 15195 2918 15204
rect 7610 15260 7918 15269
rect 7610 15258 7616 15260
rect 7672 15258 7696 15260
rect 7752 15258 7776 15260
rect 7832 15258 7856 15260
rect 7912 15258 7918 15260
rect 7672 15206 7674 15258
rect 7854 15206 7856 15258
rect 7610 15204 7616 15206
rect 7672 15204 7696 15206
rect 7752 15204 7776 15206
rect 7832 15204 7856 15206
rect 7912 15204 7918 15206
rect 7610 15195 7918 15204
rect 12610 15260 12918 15269
rect 12610 15258 12616 15260
rect 12672 15258 12696 15260
rect 12752 15258 12776 15260
rect 12832 15258 12856 15260
rect 12912 15258 12918 15260
rect 12672 15206 12674 15258
rect 12854 15206 12856 15258
rect 12610 15204 12616 15206
rect 12672 15204 12696 15206
rect 12752 15204 12776 15206
rect 12832 15204 12856 15206
rect 12912 15204 12918 15206
rect 12610 15195 12918 15204
rect 17610 15260 17918 15269
rect 17610 15258 17616 15260
rect 17672 15258 17696 15260
rect 17752 15258 17776 15260
rect 17832 15258 17856 15260
rect 17912 15258 17918 15260
rect 17672 15206 17674 15258
rect 17854 15206 17856 15258
rect 17610 15204 17616 15206
rect 17672 15204 17696 15206
rect 17752 15204 17776 15206
rect 17832 15204 17856 15206
rect 17912 15204 17918 15206
rect 17610 15195 17918 15204
rect 22610 15260 22918 15269
rect 22610 15258 22616 15260
rect 22672 15258 22696 15260
rect 22752 15258 22776 15260
rect 22832 15258 22856 15260
rect 22912 15258 22918 15260
rect 22672 15206 22674 15258
rect 22854 15206 22856 15258
rect 22610 15204 22616 15206
rect 22672 15204 22696 15206
rect 22752 15204 22776 15206
rect 22832 15204 22856 15206
rect 22912 15204 22918 15206
rect 22610 15195 22918 15204
rect 27610 15260 27918 15269
rect 27610 15258 27616 15260
rect 27672 15258 27696 15260
rect 27752 15258 27776 15260
rect 27832 15258 27856 15260
rect 27912 15258 27918 15260
rect 27672 15206 27674 15258
rect 27854 15206 27856 15258
rect 27610 15204 27616 15206
rect 27672 15204 27696 15206
rect 27752 15204 27776 15206
rect 27832 15204 27856 15206
rect 27912 15204 27918 15206
rect 27610 15195 27918 15204
rect 32610 15260 32918 15269
rect 32610 15258 32616 15260
rect 32672 15258 32696 15260
rect 32752 15258 32776 15260
rect 32832 15258 32856 15260
rect 32912 15258 32918 15260
rect 32672 15206 32674 15258
rect 32854 15206 32856 15258
rect 32610 15204 32616 15206
rect 32672 15204 32696 15206
rect 32752 15204 32776 15206
rect 32832 15204 32856 15206
rect 32912 15204 32918 15206
rect 32610 15195 32918 15204
rect 37610 15260 37918 15269
rect 37610 15258 37616 15260
rect 37672 15258 37696 15260
rect 37752 15258 37776 15260
rect 37832 15258 37856 15260
rect 37912 15258 37918 15260
rect 37672 15206 37674 15258
rect 37854 15206 37856 15258
rect 37610 15204 37616 15206
rect 37672 15204 37696 15206
rect 37752 15204 37776 15206
rect 37832 15204 37856 15206
rect 37912 15204 37918 15206
rect 37610 15195 37918 15204
rect 1950 14716 2258 14725
rect 1950 14714 1956 14716
rect 2012 14714 2036 14716
rect 2092 14714 2116 14716
rect 2172 14714 2196 14716
rect 2252 14714 2258 14716
rect 2012 14662 2014 14714
rect 2194 14662 2196 14714
rect 1950 14660 1956 14662
rect 2012 14660 2036 14662
rect 2092 14660 2116 14662
rect 2172 14660 2196 14662
rect 2252 14660 2258 14662
rect 1950 14651 2258 14660
rect 6950 14716 7258 14725
rect 6950 14714 6956 14716
rect 7012 14714 7036 14716
rect 7092 14714 7116 14716
rect 7172 14714 7196 14716
rect 7252 14714 7258 14716
rect 7012 14662 7014 14714
rect 7194 14662 7196 14714
rect 6950 14660 6956 14662
rect 7012 14660 7036 14662
rect 7092 14660 7116 14662
rect 7172 14660 7196 14662
rect 7252 14660 7258 14662
rect 6950 14651 7258 14660
rect 11950 14716 12258 14725
rect 11950 14714 11956 14716
rect 12012 14714 12036 14716
rect 12092 14714 12116 14716
rect 12172 14714 12196 14716
rect 12252 14714 12258 14716
rect 12012 14662 12014 14714
rect 12194 14662 12196 14714
rect 11950 14660 11956 14662
rect 12012 14660 12036 14662
rect 12092 14660 12116 14662
rect 12172 14660 12196 14662
rect 12252 14660 12258 14662
rect 11950 14651 12258 14660
rect 16950 14716 17258 14725
rect 16950 14714 16956 14716
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17252 14714 17258 14716
rect 17012 14662 17014 14714
rect 17194 14662 17196 14714
rect 16950 14660 16956 14662
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 17252 14660 17258 14662
rect 16950 14651 17258 14660
rect 21950 14716 22258 14725
rect 21950 14714 21956 14716
rect 22012 14714 22036 14716
rect 22092 14714 22116 14716
rect 22172 14714 22196 14716
rect 22252 14714 22258 14716
rect 22012 14662 22014 14714
rect 22194 14662 22196 14714
rect 21950 14660 21956 14662
rect 22012 14660 22036 14662
rect 22092 14660 22116 14662
rect 22172 14660 22196 14662
rect 22252 14660 22258 14662
rect 21950 14651 22258 14660
rect 26950 14716 27258 14725
rect 26950 14714 26956 14716
rect 27012 14714 27036 14716
rect 27092 14714 27116 14716
rect 27172 14714 27196 14716
rect 27252 14714 27258 14716
rect 27012 14662 27014 14714
rect 27194 14662 27196 14714
rect 26950 14660 26956 14662
rect 27012 14660 27036 14662
rect 27092 14660 27116 14662
rect 27172 14660 27196 14662
rect 27252 14660 27258 14662
rect 26950 14651 27258 14660
rect 31950 14716 32258 14725
rect 31950 14714 31956 14716
rect 32012 14714 32036 14716
rect 32092 14714 32116 14716
rect 32172 14714 32196 14716
rect 32252 14714 32258 14716
rect 32012 14662 32014 14714
rect 32194 14662 32196 14714
rect 31950 14660 31956 14662
rect 32012 14660 32036 14662
rect 32092 14660 32116 14662
rect 32172 14660 32196 14662
rect 32252 14660 32258 14662
rect 31950 14651 32258 14660
rect 36950 14716 37258 14725
rect 36950 14714 36956 14716
rect 37012 14714 37036 14716
rect 37092 14714 37116 14716
rect 37172 14714 37196 14716
rect 37252 14714 37258 14716
rect 37012 14662 37014 14714
rect 37194 14662 37196 14714
rect 36950 14660 36956 14662
rect 37012 14660 37036 14662
rect 37092 14660 37116 14662
rect 37172 14660 37196 14662
rect 37252 14660 37258 14662
rect 36950 14651 37258 14660
rect 2610 14172 2918 14181
rect 2610 14170 2616 14172
rect 2672 14170 2696 14172
rect 2752 14170 2776 14172
rect 2832 14170 2856 14172
rect 2912 14170 2918 14172
rect 2672 14118 2674 14170
rect 2854 14118 2856 14170
rect 2610 14116 2616 14118
rect 2672 14116 2696 14118
rect 2752 14116 2776 14118
rect 2832 14116 2856 14118
rect 2912 14116 2918 14118
rect 2610 14107 2918 14116
rect 7610 14172 7918 14181
rect 7610 14170 7616 14172
rect 7672 14170 7696 14172
rect 7752 14170 7776 14172
rect 7832 14170 7856 14172
rect 7912 14170 7918 14172
rect 7672 14118 7674 14170
rect 7854 14118 7856 14170
rect 7610 14116 7616 14118
rect 7672 14116 7696 14118
rect 7752 14116 7776 14118
rect 7832 14116 7856 14118
rect 7912 14116 7918 14118
rect 7610 14107 7918 14116
rect 12610 14172 12918 14181
rect 12610 14170 12616 14172
rect 12672 14170 12696 14172
rect 12752 14170 12776 14172
rect 12832 14170 12856 14172
rect 12912 14170 12918 14172
rect 12672 14118 12674 14170
rect 12854 14118 12856 14170
rect 12610 14116 12616 14118
rect 12672 14116 12696 14118
rect 12752 14116 12776 14118
rect 12832 14116 12856 14118
rect 12912 14116 12918 14118
rect 12610 14107 12918 14116
rect 17610 14172 17918 14181
rect 17610 14170 17616 14172
rect 17672 14170 17696 14172
rect 17752 14170 17776 14172
rect 17832 14170 17856 14172
rect 17912 14170 17918 14172
rect 17672 14118 17674 14170
rect 17854 14118 17856 14170
rect 17610 14116 17616 14118
rect 17672 14116 17696 14118
rect 17752 14116 17776 14118
rect 17832 14116 17856 14118
rect 17912 14116 17918 14118
rect 17610 14107 17918 14116
rect 22610 14172 22918 14181
rect 22610 14170 22616 14172
rect 22672 14170 22696 14172
rect 22752 14170 22776 14172
rect 22832 14170 22856 14172
rect 22912 14170 22918 14172
rect 22672 14118 22674 14170
rect 22854 14118 22856 14170
rect 22610 14116 22616 14118
rect 22672 14116 22696 14118
rect 22752 14116 22776 14118
rect 22832 14116 22856 14118
rect 22912 14116 22918 14118
rect 22610 14107 22918 14116
rect 27610 14172 27918 14181
rect 27610 14170 27616 14172
rect 27672 14170 27696 14172
rect 27752 14170 27776 14172
rect 27832 14170 27856 14172
rect 27912 14170 27918 14172
rect 27672 14118 27674 14170
rect 27854 14118 27856 14170
rect 27610 14116 27616 14118
rect 27672 14116 27696 14118
rect 27752 14116 27776 14118
rect 27832 14116 27856 14118
rect 27912 14116 27918 14118
rect 27610 14107 27918 14116
rect 32610 14172 32918 14181
rect 32610 14170 32616 14172
rect 32672 14170 32696 14172
rect 32752 14170 32776 14172
rect 32832 14170 32856 14172
rect 32912 14170 32918 14172
rect 32672 14118 32674 14170
rect 32854 14118 32856 14170
rect 32610 14116 32616 14118
rect 32672 14116 32696 14118
rect 32752 14116 32776 14118
rect 32832 14116 32856 14118
rect 32912 14116 32918 14118
rect 32610 14107 32918 14116
rect 37610 14172 37918 14181
rect 37610 14170 37616 14172
rect 37672 14170 37696 14172
rect 37752 14170 37776 14172
rect 37832 14170 37856 14172
rect 37912 14170 37918 14172
rect 37672 14118 37674 14170
rect 37854 14118 37856 14170
rect 37610 14116 37616 14118
rect 37672 14116 37696 14118
rect 37752 14116 37776 14118
rect 37832 14116 37856 14118
rect 37912 14116 37918 14118
rect 37610 14107 37918 14116
rect 1950 13628 2258 13637
rect 1950 13626 1956 13628
rect 2012 13626 2036 13628
rect 2092 13626 2116 13628
rect 2172 13626 2196 13628
rect 2252 13626 2258 13628
rect 2012 13574 2014 13626
rect 2194 13574 2196 13626
rect 1950 13572 1956 13574
rect 2012 13572 2036 13574
rect 2092 13572 2116 13574
rect 2172 13572 2196 13574
rect 2252 13572 2258 13574
rect 1950 13563 2258 13572
rect 6950 13628 7258 13637
rect 6950 13626 6956 13628
rect 7012 13626 7036 13628
rect 7092 13626 7116 13628
rect 7172 13626 7196 13628
rect 7252 13626 7258 13628
rect 7012 13574 7014 13626
rect 7194 13574 7196 13626
rect 6950 13572 6956 13574
rect 7012 13572 7036 13574
rect 7092 13572 7116 13574
rect 7172 13572 7196 13574
rect 7252 13572 7258 13574
rect 6950 13563 7258 13572
rect 11950 13628 12258 13637
rect 11950 13626 11956 13628
rect 12012 13626 12036 13628
rect 12092 13626 12116 13628
rect 12172 13626 12196 13628
rect 12252 13626 12258 13628
rect 12012 13574 12014 13626
rect 12194 13574 12196 13626
rect 11950 13572 11956 13574
rect 12012 13572 12036 13574
rect 12092 13572 12116 13574
rect 12172 13572 12196 13574
rect 12252 13572 12258 13574
rect 11950 13563 12258 13572
rect 16950 13628 17258 13637
rect 16950 13626 16956 13628
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17252 13626 17258 13628
rect 17012 13574 17014 13626
rect 17194 13574 17196 13626
rect 16950 13572 16956 13574
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 17252 13572 17258 13574
rect 16950 13563 17258 13572
rect 21950 13628 22258 13637
rect 21950 13626 21956 13628
rect 22012 13626 22036 13628
rect 22092 13626 22116 13628
rect 22172 13626 22196 13628
rect 22252 13626 22258 13628
rect 22012 13574 22014 13626
rect 22194 13574 22196 13626
rect 21950 13572 21956 13574
rect 22012 13572 22036 13574
rect 22092 13572 22116 13574
rect 22172 13572 22196 13574
rect 22252 13572 22258 13574
rect 21950 13563 22258 13572
rect 26950 13628 27258 13637
rect 26950 13626 26956 13628
rect 27012 13626 27036 13628
rect 27092 13626 27116 13628
rect 27172 13626 27196 13628
rect 27252 13626 27258 13628
rect 27012 13574 27014 13626
rect 27194 13574 27196 13626
rect 26950 13572 26956 13574
rect 27012 13572 27036 13574
rect 27092 13572 27116 13574
rect 27172 13572 27196 13574
rect 27252 13572 27258 13574
rect 26950 13563 27258 13572
rect 31950 13628 32258 13637
rect 31950 13626 31956 13628
rect 32012 13626 32036 13628
rect 32092 13626 32116 13628
rect 32172 13626 32196 13628
rect 32252 13626 32258 13628
rect 32012 13574 32014 13626
rect 32194 13574 32196 13626
rect 31950 13572 31956 13574
rect 32012 13572 32036 13574
rect 32092 13572 32116 13574
rect 32172 13572 32196 13574
rect 32252 13572 32258 13574
rect 31950 13563 32258 13572
rect 36950 13628 37258 13637
rect 36950 13626 36956 13628
rect 37012 13626 37036 13628
rect 37092 13626 37116 13628
rect 37172 13626 37196 13628
rect 37252 13626 37258 13628
rect 37012 13574 37014 13626
rect 37194 13574 37196 13626
rect 36950 13572 36956 13574
rect 37012 13572 37036 13574
rect 37092 13572 37116 13574
rect 37172 13572 37196 13574
rect 37252 13572 37258 13574
rect 36950 13563 37258 13572
rect 2610 13084 2918 13093
rect 2610 13082 2616 13084
rect 2672 13082 2696 13084
rect 2752 13082 2776 13084
rect 2832 13082 2856 13084
rect 2912 13082 2918 13084
rect 2672 13030 2674 13082
rect 2854 13030 2856 13082
rect 2610 13028 2616 13030
rect 2672 13028 2696 13030
rect 2752 13028 2776 13030
rect 2832 13028 2856 13030
rect 2912 13028 2918 13030
rect 2610 13019 2918 13028
rect 7610 13084 7918 13093
rect 7610 13082 7616 13084
rect 7672 13082 7696 13084
rect 7752 13082 7776 13084
rect 7832 13082 7856 13084
rect 7912 13082 7918 13084
rect 7672 13030 7674 13082
rect 7854 13030 7856 13082
rect 7610 13028 7616 13030
rect 7672 13028 7696 13030
rect 7752 13028 7776 13030
rect 7832 13028 7856 13030
rect 7912 13028 7918 13030
rect 7610 13019 7918 13028
rect 12610 13084 12918 13093
rect 12610 13082 12616 13084
rect 12672 13082 12696 13084
rect 12752 13082 12776 13084
rect 12832 13082 12856 13084
rect 12912 13082 12918 13084
rect 12672 13030 12674 13082
rect 12854 13030 12856 13082
rect 12610 13028 12616 13030
rect 12672 13028 12696 13030
rect 12752 13028 12776 13030
rect 12832 13028 12856 13030
rect 12912 13028 12918 13030
rect 12610 13019 12918 13028
rect 17610 13084 17918 13093
rect 17610 13082 17616 13084
rect 17672 13082 17696 13084
rect 17752 13082 17776 13084
rect 17832 13082 17856 13084
rect 17912 13082 17918 13084
rect 17672 13030 17674 13082
rect 17854 13030 17856 13082
rect 17610 13028 17616 13030
rect 17672 13028 17696 13030
rect 17752 13028 17776 13030
rect 17832 13028 17856 13030
rect 17912 13028 17918 13030
rect 17610 13019 17918 13028
rect 22610 13084 22918 13093
rect 22610 13082 22616 13084
rect 22672 13082 22696 13084
rect 22752 13082 22776 13084
rect 22832 13082 22856 13084
rect 22912 13082 22918 13084
rect 22672 13030 22674 13082
rect 22854 13030 22856 13082
rect 22610 13028 22616 13030
rect 22672 13028 22696 13030
rect 22752 13028 22776 13030
rect 22832 13028 22856 13030
rect 22912 13028 22918 13030
rect 22610 13019 22918 13028
rect 27610 13084 27918 13093
rect 27610 13082 27616 13084
rect 27672 13082 27696 13084
rect 27752 13082 27776 13084
rect 27832 13082 27856 13084
rect 27912 13082 27918 13084
rect 27672 13030 27674 13082
rect 27854 13030 27856 13082
rect 27610 13028 27616 13030
rect 27672 13028 27696 13030
rect 27752 13028 27776 13030
rect 27832 13028 27856 13030
rect 27912 13028 27918 13030
rect 27610 13019 27918 13028
rect 32610 13084 32918 13093
rect 32610 13082 32616 13084
rect 32672 13082 32696 13084
rect 32752 13082 32776 13084
rect 32832 13082 32856 13084
rect 32912 13082 32918 13084
rect 32672 13030 32674 13082
rect 32854 13030 32856 13082
rect 32610 13028 32616 13030
rect 32672 13028 32696 13030
rect 32752 13028 32776 13030
rect 32832 13028 32856 13030
rect 32912 13028 32918 13030
rect 32610 13019 32918 13028
rect 37610 13084 37918 13093
rect 37610 13082 37616 13084
rect 37672 13082 37696 13084
rect 37752 13082 37776 13084
rect 37832 13082 37856 13084
rect 37912 13082 37918 13084
rect 37672 13030 37674 13082
rect 37854 13030 37856 13082
rect 37610 13028 37616 13030
rect 37672 13028 37696 13030
rect 37752 13028 37776 13030
rect 37832 13028 37856 13030
rect 37912 13028 37918 13030
rect 37610 13019 37918 13028
rect 1950 12540 2258 12549
rect 1950 12538 1956 12540
rect 2012 12538 2036 12540
rect 2092 12538 2116 12540
rect 2172 12538 2196 12540
rect 2252 12538 2258 12540
rect 2012 12486 2014 12538
rect 2194 12486 2196 12538
rect 1950 12484 1956 12486
rect 2012 12484 2036 12486
rect 2092 12484 2116 12486
rect 2172 12484 2196 12486
rect 2252 12484 2258 12486
rect 1950 12475 2258 12484
rect 6950 12540 7258 12549
rect 6950 12538 6956 12540
rect 7012 12538 7036 12540
rect 7092 12538 7116 12540
rect 7172 12538 7196 12540
rect 7252 12538 7258 12540
rect 7012 12486 7014 12538
rect 7194 12486 7196 12538
rect 6950 12484 6956 12486
rect 7012 12484 7036 12486
rect 7092 12484 7116 12486
rect 7172 12484 7196 12486
rect 7252 12484 7258 12486
rect 6950 12475 7258 12484
rect 11950 12540 12258 12549
rect 11950 12538 11956 12540
rect 12012 12538 12036 12540
rect 12092 12538 12116 12540
rect 12172 12538 12196 12540
rect 12252 12538 12258 12540
rect 12012 12486 12014 12538
rect 12194 12486 12196 12538
rect 11950 12484 11956 12486
rect 12012 12484 12036 12486
rect 12092 12484 12116 12486
rect 12172 12484 12196 12486
rect 12252 12484 12258 12486
rect 11950 12475 12258 12484
rect 16950 12540 17258 12549
rect 16950 12538 16956 12540
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17252 12538 17258 12540
rect 17012 12486 17014 12538
rect 17194 12486 17196 12538
rect 16950 12484 16956 12486
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 17252 12484 17258 12486
rect 16950 12475 17258 12484
rect 21950 12540 22258 12549
rect 21950 12538 21956 12540
rect 22012 12538 22036 12540
rect 22092 12538 22116 12540
rect 22172 12538 22196 12540
rect 22252 12538 22258 12540
rect 22012 12486 22014 12538
rect 22194 12486 22196 12538
rect 21950 12484 21956 12486
rect 22012 12484 22036 12486
rect 22092 12484 22116 12486
rect 22172 12484 22196 12486
rect 22252 12484 22258 12486
rect 21950 12475 22258 12484
rect 26950 12540 27258 12549
rect 26950 12538 26956 12540
rect 27012 12538 27036 12540
rect 27092 12538 27116 12540
rect 27172 12538 27196 12540
rect 27252 12538 27258 12540
rect 27012 12486 27014 12538
rect 27194 12486 27196 12538
rect 26950 12484 26956 12486
rect 27012 12484 27036 12486
rect 27092 12484 27116 12486
rect 27172 12484 27196 12486
rect 27252 12484 27258 12486
rect 26950 12475 27258 12484
rect 31950 12540 32258 12549
rect 31950 12538 31956 12540
rect 32012 12538 32036 12540
rect 32092 12538 32116 12540
rect 32172 12538 32196 12540
rect 32252 12538 32258 12540
rect 32012 12486 32014 12538
rect 32194 12486 32196 12538
rect 31950 12484 31956 12486
rect 32012 12484 32036 12486
rect 32092 12484 32116 12486
rect 32172 12484 32196 12486
rect 32252 12484 32258 12486
rect 31950 12475 32258 12484
rect 36950 12540 37258 12549
rect 36950 12538 36956 12540
rect 37012 12538 37036 12540
rect 37092 12538 37116 12540
rect 37172 12538 37196 12540
rect 37252 12538 37258 12540
rect 37012 12486 37014 12538
rect 37194 12486 37196 12538
rect 36950 12484 36956 12486
rect 37012 12484 37036 12486
rect 37092 12484 37116 12486
rect 37172 12484 37196 12486
rect 37252 12484 37258 12486
rect 36950 12475 37258 12484
rect 2610 11996 2918 12005
rect 2610 11994 2616 11996
rect 2672 11994 2696 11996
rect 2752 11994 2776 11996
rect 2832 11994 2856 11996
rect 2912 11994 2918 11996
rect 2672 11942 2674 11994
rect 2854 11942 2856 11994
rect 2610 11940 2616 11942
rect 2672 11940 2696 11942
rect 2752 11940 2776 11942
rect 2832 11940 2856 11942
rect 2912 11940 2918 11942
rect 2610 11931 2918 11940
rect 7610 11996 7918 12005
rect 7610 11994 7616 11996
rect 7672 11994 7696 11996
rect 7752 11994 7776 11996
rect 7832 11994 7856 11996
rect 7912 11994 7918 11996
rect 7672 11942 7674 11994
rect 7854 11942 7856 11994
rect 7610 11940 7616 11942
rect 7672 11940 7696 11942
rect 7752 11940 7776 11942
rect 7832 11940 7856 11942
rect 7912 11940 7918 11942
rect 7610 11931 7918 11940
rect 12610 11996 12918 12005
rect 12610 11994 12616 11996
rect 12672 11994 12696 11996
rect 12752 11994 12776 11996
rect 12832 11994 12856 11996
rect 12912 11994 12918 11996
rect 12672 11942 12674 11994
rect 12854 11942 12856 11994
rect 12610 11940 12616 11942
rect 12672 11940 12696 11942
rect 12752 11940 12776 11942
rect 12832 11940 12856 11942
rect 12912 11940 12918 11942
rect 12610 11931 12918 11940
rect 17610 11996 17918 12005
rect 17610 11994 17616 11996
rect 17672 11994 17696 11996
rect 17752 11994 17776 11996
rect 17832 11994 17856 11996
rect 17912 11994 17918 11996
rect 17672 11942 17674 11994
rect 17854 11942 17856 11994
rect 17610 11940 17616 11942
rect 17672 11940 17696 11942
rect 17752 11940 17776 11942
rect 17832 11940 17856 11942
rect 17912 11940 17918 11942
rect 17610 11931 17918 11940
rect 22610 11996 22918 12005
rect 22610 11994 22616 11996
rect 22672 11994 22696 11996
rect 22752 11994 22776 11996
rect 22832 11994 22856 11996
rect 22912 11994 22918 11996
rect 22672 11942 22674 11994
rect 22854 11942 22856 11994
rect 22610 11940 22616 11942
rect 22672 11940 22696 11942
rect 22752 11940 22776 11942
rect 22832 11940 22856 11942
rect 22912 11940 22918 11942
rect 22610 11931 22918 11940
rect 27610 11996 27918 12005
rect 27610 11994 27616 11996
rect 27672 11994 27696 11996
rect 27752 11994 27776 11996
rect 27832 11994 27856 11996
rect 27912 11994 27918 11996
rect 27672 11942 27674 11994
rect 27854 11942 27856 11994
rect 27610 11940 27616 11942
rect 27672 11940 27696 11942
rect 27752 11940 27776 11942
rect 27832 11940 27856 11942
rect 27912 11940 27918 11942
rect 27610 11931 27918 11940
rect 32610 11996 32918 12005
rect 32610 11994 32616 11996
rect 32672 11994 32696 11996
rect 32752 11994 32776 11996
rect 32832 11994 32856 11996
rect 32912 11994 32918 11996
rect 32672 11942 32674 11994
rect 32854 11942 32856 11994
rect 32610 11940 32616 11942
rect 32672 11940 32696 11942
rect 32752 11940 32776 11942
rect 32832 11940 32856 11942
rect 32912 11940 32918 11942
rect 32610 11931 32918 11940
rect 37610 11996 37918 12005
rect 37610 11994 37616 11996
rect 37672 11994 37696 11996
rect 37752 11994 37776 11996
rect 37832 11994 37856 11996
rect 37912 11994 37918 11996
rect 37672 11942 37674 11994
rect 37854 11942 37856 11994
rect 37610 11940 37616 11942
rect 37672 11940 37696 11942
rect 37752 11940 37776 11942
rect 37832 11940 37856 11942
rect 37912 11940 37918 11942
rect 37610 11931 37918 11940
rect 1950 11452 2258 11461
rect 1950 11450 1956 11452
rect 2012 11450 2036 11452
rect 2092 11450 2116 11452
rect 2172 11450 2196 11452
rect 2252 11450 2258 11452
rect 2012 11398 2014 11450
rect 2194 11398 2196 11450
rect 1950 11396 1956 11398
rect 2012 11396 2036 11398
rect 2092 11396 2116 11398
rect 2172 11396 2196 11398
rect 2252 11396 2258 11398
rect 1950 11387 2258 11396
rect 6950 11452 7258 11461
rect 6950 11450 6956 11452
rect 7012 11450 7036 11452
rect 7092 11450 7116 11452
rect 7172 11450 7196 11452
rect 7252 11450 7258 11452
rect 7012 11398 7014 11450
rect 7194 11398 7196 11450
rect 6950 11396 6956 11398
rect 7012 11396 7036 11398
rect 7092 11396 7116 11398
rect 7172 11396 7196 11398
rect 7252 11396 7258 11398
rect 6950 11387 7258 11396
rect 11950 11452 12258 11461
rect 11950 11450 11956 11452
rect 12012 11450 12036 11452
rect 12092 11450 12116 11452
rect 12172 11450 12196 11452
rect 12252 11450 12258 11452
rect 12012 11398 12014 11450
rect 12194 11398 12196 11450
rect 11950 11396 11956 11398
rect 12012 11396 12036 11398
rect 12092 11396 12116 11398
rect 12172 11396 12196 11398
rect 12252 11396 12258 11398
rect 11950 11387 12258 11396
rect 16950 11452 17258 11461
rect 16950 11450 16956 11452
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17252 11450 17258 11452
rect 17012 11398 17014 11450
rect 17194 11398 17196 11450
rect 16950 11396 16956 11398
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 17252 11396 17258 11398
rect 16950 11387 17258 11396
rect 21950 11452 22258 11461
rect 21950 11450 21956 11452
rect 22012 11450 22036 11452
rect 22092 11450 22116 11452
rect 22172 11450 22196 11452
rect 22252 11450 22258 11452
rect 22012 11398 22014 11450
rect 22194 11398 22196 11450
rect 21950 11396 21956 11398
rect 22012 11396 22036 11398
rect 22092 11396 22116 11398
rect 22172 11396 22196 11398
rect 22252 11396 22258 11398
rect 21950 11387 22258 11396
rect 26950 11452 27258 11461
rect 26950 11450 26956 11452
rect 27012 11450 27036 11452
rect 27092 11450 27116 11452
rect 27172 11450 27196 11452
rect 27252 11450 27258 11452
rect 27012 11398 27014 11450
rect 27194 11398 27196 11450
rect 26950 11396 26956 11398
rect 27012 11396 27036 11398
rect 27092 11396 27116 11398
rect 27172 11396 27196 11398
rect 27252 11396 27258 11398
rect 26950 11387 27258 11396
rect 31950 11452 32258 11461
rect 31950 11450 31956 11452
rect 32012 11450 32036 11452
rect 32092 11450 32116 11452
rect 32172 11450 32196 11452
rect 32252 11450 32258 11452
rect 32012 11398 32014 11450
rect 32194 11398 32196 11450
rect 31950 11396 31956 11398
rect 32012 11396 32036 11398
rect 32092 11396 32116 11398
rect 32172 11396 32196 11398
rect 32252 11396 32258 11398
rect 31950 11387 32258 11396
rect 36950 11452 37258 11461
rect 36950 11450 36956 11452
rect 37012 11450 37036 11452
rect 37092 11450 37116 11452
rect 37172 11450 37196 11452
rect 37252 11450 37258 11452
rect 37012 11398 37014 11450
rect 37194 11398 37196 11450
rect 36950 11396 36956 11398
rect 37012 11396 37036 11398
rect 37092 11396 37116 11398
rect 37172 11396 37196 11398
rect 37252 11396 37258 11398
rect 36950 11387 37258 11396
rect 2610 10908 2918 10917
rect 2610 10906 2616 10908
rect 2672 10906 2696 10908
rect 2752 10906 2776 10908
rect 2832 10906 2856 10908
rect 2912 10906 2918 10908
rect 2672 10854 2674 10906
rect 2854 10854 2856 10906
rect 2610 10852 2616 10854
rect 2672 10852 2696 10854
rect 2752 10852 2776 10854
rect 2832 10852 2856 10854
rect 2912 10852 2918 10854
rect 2610 10843 2918 10852
rect 7610 10908 7918 10917
rect 7610 10906 7616 10908
rect 7672 10906 7696 10908
rect 7752 10906 7776 10908
rect 7832 10906 7856 10908
rect 7912 10906 7918 10908
rect 7672 10854 7674 10906
rect 7854 10854 7856 10906
rect 7610 10852 7616 10854
rect 7672 10852 7696 10854
rect 7752 10852 7776 10854
rect 7832 10852 7856 10854
rect 7912 10852 7918 10854
rect 7610 10843 7918 10852
rect 12610 10908 12918 10917
rect 12610 10906 12616 10908
rect 12672 10906 12696 10908
rect 12752 10906 12776 10908
rect 12832 10906 12856 10908
rect 12912 10906 12918 10908
rect 12672 10854 12674 10906
rect 12854 10854 12856 10906
rect 12610 10852 12616 10854
rect 12672 10852 12696 10854
rect 12752 10852 12776 10854
rect 12832 10852 12856 10854
rect 12912 10852 12918 10854
rect 12610 10843 12918 10852
rect 17610 10908 17918 10917
rect 17610 10906 17616 10908
rect 17672 10906 17696 10908
rect 17752 10906 17776 10908
rect 17832 10906 17856 10908
rect 17912 10906 17918 10908
rect 17672 10854 17674 10906
rect 17854 10854 17856 10906
rect 17610 10852 17616 10854
rect 17672 10852 17696 10854
rect 17752 10852 17776 10854
rect 17832 10852 17856 10854
rect 17912 10852 17918 10854
rect 17610 10843 17918 10852
rect 22610 10908 22918 10917
rect 22610 10906 22616 10908
rect 22672 10906 22696 10908
rect 22752 10906 22776 10908
rect 22832 10906 22856 10908
rect 22912 10906 22918 10908
rect 22672 10854 22674 10906
rect 22854 10854 22856 10906
rect 22610 10852 22616 10854
rect 22672 10852 22696 10854
rect 22752 10852 22776 10854
rect 22832 10852 22856 10854
rect 22912 10852 22918 10854
rect 22610 10843 22918 10852
rect 27610 10908 27918 10917
rect 27610 10906 27616 10908
rect 27672 10906 27696 10908
rect 27752 10906 27776 10908
rect 27832 10906 27856 10908
rect 27912 10906 27918 10908
rect 27672 10854 27674 10906
rect 27854 10854 27856 10906
rect 27610 10852 27616 10854
rect 27672 10852 27696 10854
rect 27752 10852 27776 10854
rect 27832 10852 27856 10854
rect 27912 10852 27918 10854
rect 27610 10843 27918 10852
rect 32610 10908 32918 10917
rect 32610 10906 32616 10908
rect 32672 10906 32696 10908
rect 32752 10906 32776 10908
rect 32832 10906 32856 10908
rect 32912 10906 32918 10908
rect 32672 10854 32674 10906
rect 32854 10854 32856 10906
rect 32610 10852 32616 10854
rect 32672 10852 32696 10854
rect 32752 10852 32776 10854
rect 32832 10852 32856 10854
rect 32912 10852 32918 10854
rect 32610 10843 32918 10852
rect 37610 10908 37918 10917
rect 37610 10906 37616 10908
rect 37672 10906 37696 10908
rect 37752 10906 37776 10908
rect 37832 10906 37856 10908
rect 37912 10906 37918 10908
rect 37672 10854 37674 10906
rect 37854 10854 37856 10906
rect 37610 10852 37616 10854
rect 37672 10852 37696 10854
rect 37752 10852 37776 10854
rect 37832 10852 37856 10854
rect 37912 10852 37918 10854
rect 37610 10843 37918 10852
rect 1950 10364 2258 10373
rect 1950 10362 1956 10364
rect 2012 10362 2036 10364
rect 2092 10362 2116 10364
rect 2172 10362 2196 10364
rect 2252 10362 2258 10364
rect 2012 10310 2014 10362
rect 2194 10310 2196 10362
rect 1950 10308 1956 10310
rect 2012 10308 2036 10310
rect 2092 10308 2116 10310
rect 2172 10308 2196 10310
rect 2252 10308 2258 10310
rect 1950 10299 2258 10308
rect 6950 10364 7258 10373
rect 6950 10362 6956 10364
rect 7012 10362 7036 10364
rect 7092 10362 7116 10364
rect 7172 10362 7196 10364
rect 7252 10362 7258 10364
rect 7012 10310 7014 10362
rect 7194 10310 7196 10362
rect 6950 10308 6956 10310
rect 7012 10308 7036 10310
rect 7092 10308 7116 10310
rect 7172 10308 7196 10310
rect 7252 10308 7258 10310
rect 6950 10299 7258 10308
rect 11950 10364 12258 10373
rect 11950 10362 11956 10364
rect 12012 10362 12036 10364
rect 12092 10362 12116 10364
rect 12172 10362 12196 10364
rect 12252 10362 12258 10364
rect 12012 10310 12014 10362
rect 12194 10310 12196 10362
rect 11950 10308 11956 10310
rect 12012 10308 12036 10310
rect 12092 10308 12116 10310
rect 12172 10308 12196 10310
rect 12252 10308 12258 10310
rect 11950 10299 12258 10308
rect 16950 10364 17258 10373
rect 16950 10362 16956 10364
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17252 10362 17258 10364
rect 17012 10310 17014 10362
rect 17194 10310 17196 10362
rect 16950 10308 16956 10310
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 17252 10308 17258 10310
rect 16950 10299 17258 10308
rect 21950 10364 22258 10373
rect 21950 10362 21956 10364
rect 22012 10362 22036 10364
rect 22092 10362 22116 10364
rect 22172 10362 22196 10364
rect 22252 10362 22258 10364
rect 22012 10310 22014 10362
rect 22194 10310 22196 10362
rect 21950 10308 21956 10310
rect 22012 10308 22036 10310
rect 22092 10308 22116 10310
rect 22172 10308 22196 10310
rect 22252 10308 22258 10310
rect 21950 10299 22258 10308
rect 26950 10364 27258 10373
rect 26950 10362 26956 10364
rect 27012 10362 27036 10364
rect 27092 10362 27116 10364
rect 27172 10362 27196 10364
rect 27252 10362 27258 10364
rect 27012 10310 27014 10362
rect 27194 10310 27196 10362
rect 26950 10308 26956 10310
rect 27012 10308 27036 10310
rect 27092 10308 27116 10310
rect 27172 10308 27196 10310
rect 27252 10308 27258 10310
rect 26950 10299 27258 10308
rect 31950 10364 32258 10373
rect 31950 10362 31956 10364
rect 32012 10362 32036 10364
rect 32092 10362 32116 10364
rect 32172 10362 32196 10364
rect 32252 10362 32258 10364
rect 32012 10310 32014 10362
rect 32194 10310 32196 10362
rect 31950 10308 31956 10310
rect 32012 10308 32036 10310
rect 32092 10308 32116 10310
rect 32172 10308 32196 10310
rect 32252 10308 32258 10310
rect 31950 10299 32258 10308
rect 36950 10364 37258 10373
rect 36950 10362 36956 10364
rect 37012 10362 37036 10364
rect 37092 10362 37116 10364
rect 37172 10362 37196 10364
rect 37252 10362 37258 10364
rect 37012 10310 37014 10362
rect 37194 10310 37196 10362
rect 36950 10308 36956 10310
rect 37012 10308 37036 10310
rect 37092 10308 37116 10310
rect 37172 10308 37196 10310
rect 37252 10308 37258 10310
rect 36950 10299 37258 10308
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 7610 9820 7918 9829
rect 7610 9818 7616 9820
rect 7672 9818 7696 9820
rect 7752 9818 7776 9820
rect 7832 9818 7856 9820
rect 7912 9818 7918 9820
rect 7672 9766 7674 9818
rect 7854 9766 7856 9818
rect 7610 9764 7616 9766
rect 7672 9764 7696 9766
rect 7752 9764 7776 9766
rect 7832 9764 7856 9766
rect 7912 9764 7918 9766
rect 7610 9755 7918 9764
rect 12610 9820 12918 9829
rect 12610 9818 12616 9820
rect 12672 9818 12696 9820
rect 12752 9818 12776 9820
rect 12832 9818 12856 9820
rect 12912 9818 12918 9820
rect 12672 9766 12674 9818
rect 12854 9766 12856 9818
rect 12610 9764 12616 9766
rect 12672 9764 12696 9766
rect 12752 9764 12776 9766
rect 12832 9764 12856 9766
rect 12912 9764 12918 9766
rect 12610 9755 12918 9764
rect 17610 9820 17918 9829
rect 17610 9818 17616 9820
rect 17672 9818 17696 9820
rect 17752 9818 17776 9820
rect 17832 9818 17856 9820
rect 17912 9818 17918 9820
rect 17672 9766 17674 9818
rect 17854 9766 17856 9818
rect 17610 9764 17616 9766
rect 17672 9764 17696 9766
rect 17752 9764 17776 9766
rect 17832 9764 17856 9766
rect 17912 9764 17918 9766
rect 17610 9755 17918 9764
rect 22610 9820 22918 9829
rect 22610 9818 22616 9820
rect 22672 9818 22696 9820
rect 22752 9818 22776 9820
rect 22832 9818 22856 9820
rect 22912 9818 22918 9820
rect 22672 9766 22674 9818
rect 22854 9766 22856 9818
rect 22610 9764 22616 9766
rect 22672 9764 22696 9766
rect 22752 9764 22776 9766
rect 22832 9764 22856 9766
rect 22912 9764 22918 9766
rect 22610 9755 22918 9764
rect 27610 9820 27918 9829
rect 27610 9818 27616 9820
rect 27672 9818 27696 9820
rect 27752 9818 27776 9820
rect 27832 9818 27856 9820
rect 27912 9818 27918 9820
rect 27672 9766 27674 9818
rect 27854 9766 27856 9818
rect 27610 9764 27616 9766
rect 27672 9764 27696 9766
rect 27752 9764 27776 9766
rect 27832 9764 27856 9766
rect 27912 9764 27918 9766
rect 27610 9755 27918 9764
rect 32610 9820 32918 9829
rect 32610 9818 32616 9820
rect 32672 9818 32696 9820
rect 32752 9818 32776 9820
rect 32832 9818 32856 9820
rect 32912 9818 32918 9820
rect 32672 9766 32674 9818
rect 32854 9766 32856 9818
rect 32610 9764 32616 9766
rect 32672 9764 32696 9766
rect 32752 9764 32776 9766
rect 32832 9764 32856 9766
rect 32912 9764 32918 9766
rect 32610 9755 32918 9764
rect 37610 9820 37918 9829
rect 37610 9818 37616 9820
rect 37672 9818 37696 9820
rect 37752 9818 37776 9820
rect 37832 9818 37856 9820
rect 37912 9818 37918 9820
rect 37672 9766 37674 9818
rect 37854 9766 37856 9818
rect 37610 9764 37616 9766
rect 37672 9764 37696 9766
rect 37752 9764 37776 9766
rect 37832 9764 37856 9766
rect 37912 9764 37918 9766
rect 37610 9755 37918 9764
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 6950 9276 7258 9285
rect 6950 9274 6956 9276
rect 7012 9274 7036 9276
rect 7092 9274 7116 9276
rect 7172 9274 7196 9276
rect 7252 9274 7258 9276
rect 7012 9222 7014 9274
rect 7194 9222 7196 9274
rect 6950 9220 6956 9222
rect 7012 9220 7036 9222
rect 7092 9220 7116 9222
rect 7172 9220 7196 9222
rect 7252 9220 7258 9222
rect 6950 9211 7258 9220
rect 11950 9276 12258 9285
rect 11950 9274 11956 9276
rect 12012 9274 12036 9276
rect 12092 9274 12116 9276
rect 12172 9274 12196 9276
rect 12252 9274 12258 9276
rect 12012 9222 12014 9274
rect 12194 9222 12196 9274
rect 11950 9220 11956 9222
rect 12012 9220 12036 9222
rect 12092 9220 12116 9222
rect 12172 9220 12196 9222
rect 12252 9220 12258 9222
rect 11950 9211 12258 9220
rect 16950 9276 17258 9285
rect 16950 9274 16956 9276
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17252 9274 17258 9276
rect 17012 9222 17014 9274
rect 17194 9222 17196 9274
rect 16950 9220 16956 9222
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 17252 9220 17258 9222
rect 16950 9211 17258 9220
rect 21950 9276 22258 9285
rect 21950 9274 21956 9276
rect 22012 9274 22036 9276
rect 22092 9274 22116 9276
rect 22172 9274 22196 9276
rect 22252 9274 22258 9276
rect 22012 9222 22014 9274
rect 22194 9222 22196 9274
rect 21950 9220 21956 9222
rect 22012 9220 22036 9222
rect 22092 9220 22116 9222
rect 22172 9220 22196 9222
rect 22252 9220 22258 9222
rect 21950 9211 22258 9220
rect 26950 9276 27258 9285
rect 26950 9274 26956 9276
rect 27012 9274 27036 9276
rect 27092 9274 27116 9276
rect 27172 9274 27196 9276
rect 27252 9274 27258 9276
rect 27012 9222 27014 9274
rect 27194 9222 27196 9274
rect 26950 9220 26956 9222
rect 27012 9220 27036 9222
rect 27092 9220 27116 9222
rect 27172 9220 27196 9222
rect 27252 9220 27258 9222
rect 26950 9211 27258 9220
rect 31950 9276 32258 9285
rect 31950 9274 31956 9276
rect 32012 9274 32036 9276
rect 32092 9274 32116 9276
rect 32172 9274 32196 9276
rect 32252 9274 32258 9276
rect 32012 9222 32014 9274
rect 32194 9222 32196 9274
rect 31950 9220 31956 9222
rect 32012 9220 32036 9222
rect 32092 9220 32116 9222
rect 32172 9220 32196 9222
rect 32252 9220 32258 9222
rect 31950 9211 32258 9220
rect 36950 9276 37258 9285
rect 36950 9274 36956 9276
rect 37012 9274 37036 9276
rect 37092 9274 37116 9276
rect 37172 9274 37196 9276
rect 37252 9274 37258 9276
rect 37012 9222 37014 9274
rect 37194 9222 37196 9274
rect 36950 9220 36956 9222
rect 37012 9220 37036 9222
rect 37092 9220 37116 9222
rect 37172 9220 37196 9222
rect 37252 9220 37258 9222
rect 36950 9211 37258 9220
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 7610 8732 7918 8741
rect 7610 8730 7616 8732
rect 7672 8730 7696 8732
rect 7752 8730 7776 8732
rect 7832 8730 7856 8732
rect 7912 8730 7918 8732
rect 7672 8678 7674 8730
rect 7854 8678 7856 8730
rect 7610 8676 7616 8678
rect 7672 8676 7696 8678
rect 7752 8676 7776 8678
rect 7832 8676 7856 8678
rect 7912 8676 7918 8678
rect 7610 8667 7918 8676
rect 12610 8732 12918 8741
rect 12610 8730 12616 8732
rect 12672 8730 12696 8732
rect 12752 8730 12776 8732
rect 12832 8730 12856 8732
rect 12912 8730 12918 8732
rect 12672 8678 12674 8730
rect 12854 8678 12856 8730
rect 12610 8676 12616 8678
rect 12672 8676 12696 8678
rect 12752 8676 12776 8678
rect 12832 8676 12856 8678
rect 12912 8676 12918 8678
rect 12610 8667 12918 8676
rect 17610 8732 17918 8741
rect 17610 8730 17616 8732
rect 17672 8730 17696 8732
rect 17752 8730 17776 8732
rect 17832 8730 17856 8732
rect 17912 8730 17918 8732
rect 17672 8678 17674 8730
rect 17854 8678 17856 8730
rect 17610 8676 17616 8678
rect 17672 8676 17696 8678
rect 17752 8676 17776 8678
rect 17832 8676 17856 8678
rect 17912 8676 17918 8678
rect 17610 8667 17918 8676
rect 22610 8732 22918 8741
rect 22610 8730 22616 8732
rect 22672 8730 22696 8732
rect 22752 8730 22776 8732
rect 22832 8730 22856 8732
rect 22912 8730 22918 8732
rect 22672 8678 22674 8730
rect 22854 8678 22856 8730
rect 22610 8676 22616 8678
rect 22672 8676 22696 8678
rect 22752 8676 22776 8678
rect 22832 8676 22856 8678
rect 22912 8676 22918 8678
rect 22610 8667 22918 8676
rect 27610 8732 27918 8741
rect 27610 8730 27616 8732
rect 27672 8730 27696 8732
rect 27752 8730 27776 8732
rect 27832 8730 27856 8732
rect 27912 8730 27918 8732
rect 27672 8678 27674 8730
rect 27854 8678 27856 8730
rect 27610 8676 27616 8678
rect 27672 8676 27696 8678
rect 27752 8676 27776 8678
rect 27832 8676 27856 8678
rect 27912 8676 27918 8678
rect 27610 8667 27918 8676
rect 32610 8732 32918 8741
rect 32610 8730 32616 8732
rect 32672 8730 32696 8732
rect 32752 8730 32776 8732
rect 32832 8730 32856 8732
rect 32912 8730 32918 8732
rect 32672 8678 32674 8730
rect 32854 8678 32856 8730
rect 32610 8676 32616 8678
rect 32672 8676 32696 8678
rect 32752 8676 32776 8678
rect 32832 8676 32856 8678
rect 32912 8676 32918 8678
rect 32610 8667 32918 8676
rect 37610 8732 37918 8741
rect 37610 8730 37616 8732
rect 37672 8730 37696 8732
rect 37752 8730 37776 8732
rect 37832 8730 37856 8732
rect 37912 8730 37918 8732
rect 37672 8678 37674 8730
rect 37854 8678 37856 8730
rect 37610 8676 37616 8678
rect 37672 8676 37696 8678
rect 37752 8676 37776 8678
rect 37832 8676 37856 8678
rect 37912 8676 37918 8678
rect 37610 8667 37918 8676
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 6950 8188 7258 8197
rect 6950 8186 6956 8188
rect 7012 8186 7036 8188
rect 7092 8186 7116 8188
rect 7172 8186 7196 8188
rect 7252 8186 7258 8188
rect 7012 8134 7014 8186
rect 7194 8134 7196 8186
rect 6950 8132 6956 8134
rect 7012 8132 7036 8134
rect 7092 8132 7116 8134
rect 7172 8132 7196 8134
rect 7252 8132 7258 8134
rect 6950 8123 7258 8132
rect 11950 8188 12258 8197
rect 11950 8186 11956 8188
rect 12012 8186 12036 8188
rect 12092 8186 12116 8188
rect 12172 8186 12196 8188
rect 12252 8186 12258 8188
rect 12012 8134 12014 8186
rect 12194 8134 12196 8186
rect 11950 8132 11956 8134
rect 12012 8132 12036 8134
rect 12092 8132 12116 8134
rect 12172 8132 12196 8134
rect 12252 8132 12258 8134
rect 11950 8123 12258 8132
rect 16950 8188 17258 8197
rect 16950 8186 16956 8188
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17252 8186 17258 8188
rect 17012 8134 17014 8186
rect 17194 8134 17196 8186
rect 16950 8132 16956 8134
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 17252 8132 17258 8134
rect 16950 8123 17258 8132
rect 21950 8188 22258 8197
rect 21950 8186 21956 8188
rect 22012 8186 22036 8188
rect 22092 8186 22116 8188
rect 22172 8186 22196 8188
rect 22252 8186 22258 8188
rect 22012 8134 22014 8186
rect 22194 8134 22196 8186
rect 21950 8132 21956 8134
rect 22012 8132 22036 8134
rect 22092 8132 22116 8134
rect 22172 8132 22196 8134
rect 22252 8132 22258 8134
rect 21950 8123 22258 8132
rect 26950 8188 27258 8197
rect 26950 8186 26956 8188
rect 27012 8186 27036 8188
rect 27092 8186 27116 8188
rect 27172 8186 27196 8188
rect 27252 8186 27258 8188
rect 27012 8134 27014 8186
rect 27194 8134 27196 8186
rect 26950 8132 26956 8134
rect 27012 8132 27036 8134
rect 27092 8132 27116 8134
rect 27172 8132 27196 8134
rect 27252 8132 27258 8134
rect 26950 8123 27258 8132
rect 31950 8188 32258 8197
rect 31950 8186 31956 8188
rect 32012 8186 32036 8188
rect 32092 8186 32116 8188
rect 32172 8186 32196 8188
rect 32252 8186 32258 8188
rect 32012 8134 32014 8186
rect 32194 8134 32196 8186
rect 31950 8132 31956 8134
rect 32012 8132 32036 8134
rect 32092 8132 32116 8134
rect 32172 8132 32196 8134
rect 32252 8132 32258 8134
rect 31950 8123 32258 8132
rect 36950 8188 37258 8197
rect 36950 8186 36956 8188
rect 37012 8186 37036 8188
rect 37092 8186 37116 8188
rect 37172 8186 37196 8188
rect 37252 8186 37258 8188
rect 37012 8134 37014 8186
rect 37194 8134 37196 8186
rect 36950 8132 36956 8134
rect 37012 8132 37036 8134
rect 37092 8132 37116 8134
rect 37172 8132 37196 8134
rect 37252 8132 37258 8134
rect 36950 8123 37258 8132
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 7610 7644 7918 7653
rect 7610 7642 7616 7644
rect 7672 7642 7696 7644
rect 7752 7642 7776 7644
rect 7832 7642 7856 7644
rect 7912 7642 7918 7644
rect 7672 7590 7674 7642
rect 7854 7590 7856 7642
rect 7610 7588 7616 7590
rect 7672 7588 7696 7590
rect 7752 7588 7776 7590
rect 7832 7588 7856 7590
rect 7912 7588 7918 7590
rect 7610 7579 7918 7588
rect 12610 7644 12918 7653
rect 12610 7642 12616 7644
rect 12672 7642 12696 7644
rect 12752 7642 12776 7644
rect 12832 7642 12856 7644
rect 12912 7642 12918 7644
rect 12672 7590 12674 7642
rect 12854 7590 12856 7642
rect 12610 7588 12616 7590
rect 12672 7588 12696 7590
rect 12752 7588 12776 7590
rect 12832 7588 12856 7590
rect 12912 7588 12918 7590
rect 12610 7579 12918 7588
rect 17610 7644 17918 7653
rect 17610 7642 17616 7644
rect 17672 7642 17696 7644
rect 17752 7642 17776 7644
rect 17832 7642 17856 7644
rect 17912 7642 17918 7644
rect 17672 7590 17674 7642
rect 17854 7590 17856 7642
rect 17610 7588 17616 7590
rect 17672 7588 17696 7590
rect 17752 7588 17776 7590
rect 17832 7588 17856 7590
rect 17912 7588 17918 7590
rect 17610 7579 17918 7588
rect 22610 7644 22918 7653
rect 22610 7642 22616 7644
rect 22672 7642 22696 7644
rect 22752 7642 22776 7644
rect 22832 7642 22856 7644
rect 22912 7642 22918 7644
rect 22672 7590 22674 7642
rect 22854 7590 22856 7642
rect 22610 7588 22616 7590
rect 22672 7588 22696 7590
rect 22752 7588 22776 7590
rect 22832 7588 22856 7590
rect 22912 7588 22918 7590
rect 22610 7579 22918 7588
rect 27610 7644 27918 7653
rect 27610 7642 27616 7644
rect 27672 7642 27696 7644
rect 27752 7642 27776 7644
rect 27832 7642 27856 7644
rect 27912 7642 27918 7644
rect 27672 7590 27674 7642
rect 27854 7590 27856 7642
rect 27610 7588 27616 7590
rect 27672 7588 27696 7590
rect 27752 7588 27776 7590
rect 27832 7588 27856 7590
rect 27912 7588 27918 7590
rect 27610 7579 27918 7588
rect 32610 7644 32918 7653
rect 32610 7642 32616 7644
rect 32672 7642 32696 7644
rect 32752 7642 32776 7644
rect 32832 7642 32856 7644
rect 32912 7642 32918 7644
rect 32672 7590 32674 7642
rect 32854 7590 32856 7642
rect 32610 7588 32616 7590
rect 32672 7588 32696 7590
rect 32752 7588 32776 7590
rect 32832 7588 32856 7590
rect 32912 7588 32918 7590
rect 32610 7579 32918 7588
rect 37610 7644 37918 7653
rect 37610 7642 37616 7644
rect 37672 7642 37696 7644
rect 37752 7642 37776 7644
rect 37832 7642 37856 7644
rect 37912 7642 37918 7644
rect 37672 7590 37674 7642
rect 37854 7590 37856 7642
rect 37610 7588 37616 7590
rect 37672 7588 37696 7590
rect 37752 7588 37776 7590
rect 37832 7588 37856 7590
rect 37912 7588 37918 7590
rect 37610 7579 37918 7588
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 6950 7100 7258 7109
rect 6950 7098 6956 7100
rect 7012 7098 7036 7100
rect 7092 7098 7116 7100
rect 7172 7098 7196 7100
rect 7252 7098 7258 7100
rect 7012 7046 7014 7098
rect 7194 7046 7196 7098
rect 6950 7044 6956 7046
rect 7012 7044 7036 7046
rect 7092 7044 7116 7046
rect 7172 7044 7196 7046
rect 7252 7044 7258 7046
rect 6950 7035 7258 7044
rect 11950 7100 12258 7109
rect 11950 7098 11956 7100
rect 12012 7098 12036 7100
rect 12092 7098 12116 7100
rect 12172 7098 12196 7100
rect 12252 7098 12258 7100
rect 12012 7046 12014 7098
rect 12194 7046 12196 7098
rect 11950 7044 11956 7046
rect 12012 7044 12036 7046
rect 12092 7044 12116 7046
rect 12172 7044 12196 7046
rect 12252 7044 12258 7046
rect 11950 7035 12258 7044
rect 16950 7100 17258 7109
rect 16950 7098 16956 7100
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17252 7098 17258 7100
rect 17012 7046 17014 7098
rect 17194 7046 17196 7098
rect 16950 7044 16956 7046
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 17252 7044 17258 7046
rect 16950 7035 17258 7044
rect 21950 7100 22258 7109
rect 21950 7098 21956 7100
rect 22012 7098 22036 7100
rect 22092 7098 22116 7100
rect 22172 7098 22196 7100
rect 22252 7098 22258 7100
rect 22012 7046 22014 7098
rect 22194 7046 22196 7098
rect 21950 7044 21956 7046
rect 22012 7044 22036 7046
rect 22092 7044 22116 7046
rect 22172 7044 22196 7046
rect 22252 7044 22258 7046
rect 21950 7035 22258 7044
rect 26950 7100 27258 7109
rect 26950 7098 26956 7100
rect 27012 7098 27036 7100
rect 27092 7098 27116 7100
rect 27172 7098 27196 7100
rect 27252 7098 27258 7100
rect 27012 7046 27014 7098
rect 27194 7046 27196 7098
rect 26950 7044 26956 7046
rect 27012 7044 27036 7046
rect 27092 7044 27116 7046
rect 27172 7044 27196 7046
rect 27252 7044 27258 7046
rect 26950 7035 27258 7044
rect 31950 7100 32258 7109
rect 31950 7098 31956 7100
rect 32012 7098 32036 7100
rect 32092 7098 32116 7100
rect 32172 7098 32196 7100
rect 32252 7098 32258 7100
rect 32012 7046 32014 7098
rect 32194 7046 32196 7098
rect 31950 7044 31956 7046
rect 32012 7044 32036 7046
rect 32092 7044 32116 7046
rect 32172 7044 32196 7046
rect 32252 7044 32258 7046
rect 31950 7035 32258 7044
rect 36950 7100 37258 7109
rect 36950 7098 36956 7100
rect 37012 7098 37036 7100
rect 37092 7098 37116 7100
rect 37172 7098 37196 7100
rect 37252 7098 37258 7100
rect 37012 7046 37014 7098
rect 37194 7046 37196 7098
rect 36950 7044 36956 7046
rect 37012 7044 37036 7046
rect 37092 7044 37116 7046
rect 37172 7044 37196 7046
rect 37252 7044 37258 7046
rect 36950 7035 37258 7044
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 7610 6556 7918 6565
rect 7610 6554 7616 6556
rect 7672 6554 7696 6556
rect 7752 6554 7776 6556
rect 7832 6554 7856 6556
rect 7912 6554 7918 6556
rect 7672 6502 7674 6554
rect 7854 6502 7856 6554
rect 7610 6500 7616 6502
rect 7672 6500 7696 6502
rect 7752 6500 7776 6502
rect 7832 6500 7856 6502
rect 7912 6500 7918 6502
rect 7610 6491 7918 6500
rect 12610 6556 12918 6565
rect 12610 6554 12616 6556
rect 12672 6554 12696 6556
rect 12752 6554 12776 6556
rect 12832 6554 12856 6556
rect 12912 6554 12918 6556
rect 12672 6502 12674 6554
rect 12854 6502 12856 6554
rect 12610 6500 12616 6502
rect 12672 6500 12696 6502
rect 12752 6500 12776 6502
rect 12832 6500 12856 6502
rect 12912 6500 12918 6502
rect 12610 6491 12918 6500
rect 17610 6556 17918 6565
rect 17610 6554 17616 6556
rect 17672 6554 17696 6556
rect 17752 6554 17776 6556
rect 17832 6554 17856 6556
rect 17912 6554 17918 6556
rect 17672 6502 17674 6554
rect 17854 6502 17856 6554
rect 17610 6500 17616 6502
rect 17672 6500 17696 6502
rect 17752 6500 17776 6502
rect 17832 6500 17856 6502
rect 17912 6500 17918 6502
rect 17610 6491 17918 6500
rect 22610 6556 22918 6565
rect 22610 6554 22616 6556
rect 22672 6554 22696 6556
rect 22752 6554 22776 6556
rect 22832 6554 22856 6556
rect 22912 6554 22918 6556
rect 22672 6502 22674 6554
rect 22854 6502 22856 6554
rect 22610 6500 22616 6502
rect 22672 6500 22696 6502
rect 22752 6500 22776 6502
rect 22832 6500 22856 6502
rect 22912 6500 22918 6502
rect 22610 6491 22918 6500
rect 27610 6556 27918 6565
rect 27610 6554 27616 6556
rect 27672 6554 27696 6556
rect 27752 6554 27776 6556
rect 27832 6554 27856 6556
rect 27912 6554 27918 6556
rect 27672 6502 27674 6554
rect 27854 6502 27856 6554
rect 27610 6500 27616 6502
rect 27672 6500 27696 6502
rect 27752 6500 27776 6502
rect 27832 6500 27856 6502
rect 27912 6500 27918 6502
rect 27610 6491 27918 6500
rect 32610 6556 32918 6565
rect 32610 6554 32616 6556
rect 32672 6554 32696 6556
rect 32752 6554 32776 6556
rect 32832 6554 32856 6556
rect 32912 6554 32918 6556
rect 32672 6502 32674 6554
rect 32854 6502 32856 6554
rect 32610 6500 32616 6502
rect 32672 6500 32696 6502
rect 32752 6500 32776 6502
rect 32832 6500 32856 6502
rect 32912 6500 32918 6502
rect 32610 6491 32918 6500
rect 37610 6556 37918 6565
rect 37610 6554 37616 6556
rect 37672 6554 37696 6556
rect 37752 6554 37776 6556
rect 37832 6554 37856 6556
rect 37912 6554 37918 6556
rect 37672 6502 37674 6554
rect 37854 6502 37856 6554
rect 37610 6500 37616 6502
rect 37672 6500 37696 6502
rect 37752 6500 37776 6502
rect 37832 6500 37856 6502
rect 37912 6500 37918 6502
rect 37610 6491 37918 6500
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 6950 6012 7258 6021
rect 6950 6010 6956 6012
rect 7012 6010 7036 6012
rect 7092 6010 7116 6012
rect 7172 6010 7196 6012
rect 7252 6010 7258 6012
rect 7012 5958 7014 6010
rect 7194 5958 7196 6010
rect 6950 5956 6956 5958
rect 7012 5956 7036 5958
rect 7092 5956 7116 5958
rect 7172 5956 7196 5958
rect 7252 5956 7258 5958
rect 6950 5947 7258 5956
rect 11950 6012 12258 6021
rect 11950 6010 11956 6012
rect 12012 6010 12036 6012
rect 12092 6010 12116 6012
rect 12172 6010 12196 6012
rect 12252 6010 12258 6012
rect 12012 5958 12014 6010
rect 12194 5958 12196 6010
rect 11950 5956 11956 5958
rect 12012 5956 12036 5958
rect 12092 5956 12116 5958
rect 12172 5956 12196 5958
rect 12252 5956 12258 5958
rect 11950 5947 12258 5956
rect 16950 6012 17258 6021
rect 16950 6010 16956 6012
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17252 6010 17258 6012
rect 17012 5958 17014 6010
rect 17194 5958 17196 6010
rect 16950 5956 16956 5958
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 17252 5956 17258 5958
rect 16950 5947 17258 5956
rect 21950 6012 22258 6021
rect 21950 6010 21956 6012
rect 22012 6010 22036 6012
rect 22092 6010 22116 6012
rect 22172 6010 22196 6012
rect 22252 6010 22258 6012
rect 22012 5958 22014 6010
rect 22194 5958 22196 6010
rect 21950 5956 21956 5958
rect 22012 5956 22036 5958
rect 22092 5956 22116 5958
rect 22172 5956 22196 5958
rect 22252 5956 22258 5958
rect 21950 5947 22258 5956
rect 26950 6012 27258 6021
rect 26950 6010 26956 6012
rect 27012 6010 27036 6012
rect 27092 6010 27116 6012
rect 27172 6010 27196 6012
rect 27252 6010 27258 6012
rect 27012 5958 27014 6010
rect 27194 5958 27196 6010
rect 26950 5956 26956 5958
rect 27012 5956 27036 5958
rect 27092 5956 27116 5958
rect 27172 5956 27196 5958
rect 27252 5956 27258 5958
rect 26950 5947 27258 5956
rect 31950 6012 32258 6021
rect 31950 6010 31956 6012
rect 32012 6010 32036 6012
rect 32092 6010 32116 6012
rect 32172 6010 32196 6012
rect 32252 6010 32258 6012
rect 32012 5958 32014 6010
rect 32194 5958 32196 6010
rect 31950 5956 31956 5958
rect 32012 5956 32036 5958
rect 32092 5956 32116 5958
rect 32172 5956 32196 5958
rect 32252 5956 32258 5958
rect 31950 5947 32258 5956
rect 36950 6012 37258 6021
rect 36950 6010 36956 6012
rect 37012 6010 37036 6012
rect 37092 6010 37116 6012
rect 37172 6010 37196 6012
rect 37252 6010 37258 6012
rect 37012 5958 37014 6010
rect 37194 5958 37196 6010
rect 36950 5956 36956 5958
rect 37012 5956 37036 5958
rect 37092 5956 37116 5958
rect 37172 5956 37196 5958
rect 37252 5956 37258 5958
rect 36950 5947 37258 5956
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 7610 5468 7918 5477
rect 7610 5466 7616 5468
rect 7672 5466 7696 5468
rect 7752 5466 7776 5468
rect 7832 5466 7856 5468
rect 7912 5466 7918 5468
rect 7672 5414 7674 5466
rect 7854 5414 7856 5466
rect 7610 5412 7616 5414
rect 7672 5412 7696 5414
rect 7752 5412 7776 5414
rect 7832 5412 7856 5414
rect 7912 5412 7918 5414
rect 7610 5403 7918 5412
rect 12610 5468 12918 5477
rect 12610 5466 12616 5468
rect 12672 5466 12696 5468
rect 12752 5466 12776 5468
rect 12832 5466 12856 5468
rect 12912 5466 12918 5468
rect 12672 5414 12674 5466
rect 12854 5414 12856 5466
rect 12610 5412 12616 5414
rect 12672 5412 12696 5414
rect 12752 5412 12776 5414
rect 12832 5412 12856 5414
rect 12912 5412 12918 5414
rect 12610 5403 12918 5412
rect 17610 5468 17918 5477
rect 17610 5466 17616 5468
rect 17672 5466 17696 5468
rect 17752 5466 17776 5468
rect 17832 5466 17856 5468
rect 17912 5466 17918 5468
rect 17672 5414 17674 5466
rect 17854 5414 17856 5466
rect 17610 5412 17616 5414
rect 17672 5412 17696 5414
rect 17752 5412 17776 5414
rect 17832 5412 17856 5414
rect 17912 5412 17918 5414
rect 17610 5403 17918 5412
rect 22610 5468 22918 5477
rect 22610 5466 22616 5468
rect 22672 5466 22696 5468
rect 22752 5466 22776 5468
rect 22832 5466 22856 5468
rect 22912 5466 22918 5468
rect 22672 5414 22674 5466
rect 22854 5414 22856 5466
rect 22610 5412 22616 5414
rect 22672 5412 22696 5414
rect 22752 5412 22776 5414
rect 22832 5412 22856 5414
rect 22912 5412 22918 5414
rect 22610 5403 22918 5412
rect 27610 5468 27918 5477
rect 27610 5466 27616 5468
rect 27672 5466 27696 5468
rect 27752 5466 27776 5468
rect 27832 5466 27856 5468
rect 27912 5466 27918 5468
rect 27672 5414 27674 5466
rect 27854 5414 27856 5466
rect 27610 5412 27616 5414
rect 27672 5412 27696 5414
rect 27752 5412 27776 5414
rect 27832 5412 27856 5414
rect 27912 5412 27918 5414
rect 27610 5403 27918 5412
rect 32610 5468 32918 5477
rect 32610 5466 32616 5468
rect 32672 5466 32696 5468
rect 32752 5466 32776 5468
rect 32832 5466 32856 5468
rect 32912 5466 32918 5468
rect 32672 5414 32674 5466
rect 32854 5414 32856 5466
rect 32610 5412 32616 5414
rect 32672 5412 32696 5414
rect 32752 5412 32776 5414
rect 32832 5412 32856 5414
rect 32912 5412 32918 5414
rect 32610 5403 32918 5412
rect 37610 5468 37918 5477
rect 37610 5466 37616 5468
rect 37672 5466 37696 5468
rect 37752 5466 37776 5468
rect 37832 5466 37856 5468
rect 37912 5466 37918 5468
rect 37672 5414 37674 5466
rect 37854 5414 37856 5466
rect 37610 5412 37616 5414
rect 37672 5412 37696 5414
rect 37752 5412 37776 5414
rect 37832 5412 37856 5414
rect 37912 5412 37918 5414
rect 37610 5403 37918 5412
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 6950 4924 7258 4933
rect 6950 4922 6956 4924
rect 7012 4922 7036 4924
rect 7092 4922 7116 4924
rect 7172 4922 7196 4924
rect 7252 4922 7258 4924
rect 7012 4870 7014 4922
rect 7194 4870 7196 4922
rect 6950 4868 6956 4870
rect 7012 4868 7036 4870
rect 7092 4868 7116 4870
rect 7172 4868 7196 4870
rect 7252 4868 7258 4870
rect 6950 4859 7258 4868
rect 11950 4924 12258 4933
rect 11950 4922 11956 4924
rect 12012 4922 12036 4924
rect 12092 4922 12116 4924
rect 12172 4922 12196 4924
rect 12252 4922 12258 4924
rect 12012 4870 12014 4922
rect 12194 4870 12196 4922
rect 11950 4868 11956 4870
rect 12012 4868 12036 4870
rect 12092 4868 12116 4870
rect 12172 4868 12196 4870
rect 12252 4868 12258 4870
rect 11950 4859 12258 4868
rect 16950 4924 17258 4933
rect 16950 4922 16956 4924
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17252 4922 17258 4924
rect 17012 4870 17014 4922
rect 17194 4870 17196 4922
rect 16950 4868 16956 4870
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 17252 4868 17258 4870
rect 16950 4859 17258 4868
rect 21950 4924 22258 4933
rect 21950 4922 21956 4924
rect 22012 4922 22036 4924
rect 22092 4922 22116 4924
rect 22172 4922 22196 4924
rect 22252 4922 22258 4924
rect 22012 4870 22014 4922
rect 22194 4870 22196 4922
rect 21950 4868 21956 4870
rect 22012 4868 22036 4870
rect 22092 4868 22116 4870
rect 22172 4868 22196 4870
rect 22252 4868 22258 4870
rect 21950 4859 22258 4868
rect 26950 4924 27258 4933
rect 26950 4922 26956 4924
rect 27012 4922 27036 4924
rect 27092 4922 27116 4924
rect 27172 4922 27196 4924
rect 27252 4922 27258 4924
rect 27012 4870 27014 4922
rect 27194 4870 27196 4922
rect 26950 4868 26956 4870
rect 27012 4868 27036 4870
rect 27092 4868 27116 4870
rect 27172 4868 27196 4870
rect 27252 4868 27258 4870
rect 26950 4859 27258 4868
rect 31950 4924 32258 4933
rect 31950 4922 31956 4924
rect 32012 4922 32036 4924
rect 32092 4922 32116 4924
rect 32172 4922 32196 4924
rect 32252 4922 32258 4924
rect 32012 4870 32014 4922
rect 32194 4870 32196 4922
rect 31950 4868 31956 4870
rect 32012 4868 32036 4870
rect 32092 4868 32116 4870
rect 32172 4868 32196 4870
rect 32252 4868 32258 4870
rect 31950 4859 32258 4868
rect 36950 4924 37258 4933
rect 36950 4922 36956 4924
rect 37012 4922 37036 4924
rect 37092 4922 37116 4924
rect 37172 4922 37196 4924
rect 37252 4922 37258 4924
rect 37012 4870 37014 4922
rect 37194 4870 37196 4922
rect 36950 4868 36956 4870
rect 37012 4868 37036 4870
rect 37092 4868 37116 4870
rect 37172 4868 37196 4870
rect 37252 4868 37258 4870
rect 36950 4859 37258 4868
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 7610 4380 7918 4389
rect 7610 4378 7616 4380
rect 7672 4378 7696 4380
rect 7752 4378 7776 4380
rect 7832 4378 7856 4380
rect 7912 4378 7918 4380
rect 7672 4326 7674 4378
rect 7854 4326 7856 4378
rect 7610 4324 7616 4326
rect 7672 4324 7696 4326
rect 7752 4324 7776 4326
rect 7832 4324 7856 4326
rect 7912 4324 7918 4326
rect 7610 4315 7918 4324
rect 12610 4380 12918 4389
rect 12610 4378 12616 4380
rect 12672 4378 12696 4380
rect 12752 4378 12776 4380
rect 12832 4378 12856 4380
rect 12912 4378 12918 4380
rect 12672 4326 12674 4378
rect 12854 4326 12856 4378
rect 12610 4324 12616 4326
rect 12672 4324 12696 4326
rect 12752 4324 12776 4326
rect 12832 4324 12856 4326
rect 12912 4324 12918 4326
rect 12610 4315 12918 4324
rect 17610 4380 17918 4389
rect 17610 4378 17616 4380
rect 17672 4378 17696 4380
rect 17752 4378 17776 4380
rect 17832 4378 17856 4380
rect 17912 4378 17918 4380
rect 17672 4326 17674 4378
rect 17854 4326 17856 4378
rect 17610 4324 17616 4326
rect 17672 4324 17696 4326
rect 17752 4324 17776 4326
rect 17832 4324 17856 4326
rect 17912 4324 17918 4326
rect 17610 4315 17918 4324
rect 22610 4380 22918 4389
rect 22610 4378 22616 4380
rect 22672 4378 22696 4380
rect 22752 4378 22776 4380
rect 22832 4378 22856 4380
rect 22912 4378 22918 4380
rect 22672 4326 22674 4378
rect 22854 4326 22856 4378
rect 22610 4324 22616 4326
rect 22672 4324 22696 4326
rect 22752 4324 22776 4326
rect 22832 4324 22856 4326
rect 22912 4324 22918 4326
rect 22610 4315 22918 4324
rect 27610 4380 27918 4389
rect 27610 4378 27616 4380
rect 27672 4378 27696 4380
rect 27752 4378 27776 4380
rect 27832 4378 27856 4380
rect 27912 4378 27918 4380
rect 27672 4326 27674 4378
rect 27854 4326 27856 4378
rect 27610 4324 27616 4326
rect 27672 4324 27696 4326
rect 27752 4324 27776 4326
rect 27832 4324 27856 4326
rect 27912 4324 27918 4326
rect 27610 4315 27918 4324
rect 32610 4380 32918 4389
rect 32610 4378 32616 4380
rect 32672 4378 32696 4380
rect 32752 4378 32776 4380
rect 32832 4378 32856 4380
rect 32912 4378 32918 4380
rect 32672 4326 32674 4378
rect 32854 4326 32856 4378
rect 32610 4324 32616 4326
rect 32672 4324 32696 4326
rect 32752 4324 32776 4326
rect 32832 4324 32856 4326
rect 32912 4324 32918 4326
rect 32610 4315 32918 4324
rect 37610 4380 37918 4389
rect 37610 4378 37616 4380
rect 37672 4378 37696 4380
rect 37752 4378 37776 4380
rect 37832 4378 37856 4380
rect 37912 4378 37918 4380
rect 37672 4326 37674 4378
rect 37854 4326 37856 4378
rect 37610 4324 37616 4326
rect 37672 4324 37696 4326
rect 37752 4324 37776 4326
rect 37832 4324 37856 4326
rect 37912 4324 37918 4326
rect 37610 4315 37918 4324
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 6950 3836 7258 3845
rect 6950 3834 6956 3836
rect 7012 3834 7036 3836
rect 7092 3834 7116 3836
rect 7172 3834 7196 3836
rect 7252 3834 7258 3836
rect 7012 3782 7014 3834
rect 7194 3782 7196 3834
rect 6950 3780 6956 3782
rect 7012 3780 7036 3782
rect 7092 3780 7116 3782
rect 7172 3780 7196 3782
rect 7252 3780 7258 3782
rect 6950 3771 7258 3780
rect 11950 3836 12258 3845
rect 11950 3834 11956 3836
rect 12012 3834 12036 3836
rect 12092 3834 12116 3836
rect 12172 3834 12196 3836
rect 12252 3834 12258 3836
rect 12012 3782 12014 3834
rect 12194 3782 12196 3834
rect 11950 3780 11956 3782
rect 12012 3780 12036 3782
rect 12092 3780 12116 3782
rect 12172 3780 12196 3782
rect 12252 3780 12258 3782
rect 11950 3771 12258 3780
rect 16950 3836 17258 3845
rect 16950 3834 16956 3836
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17252 3834 17258 3836
rect 17012 3782 17014 3834
rect 17194 3782 17196 3834
rect 16950 3780 16956 3782
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 17252 3780 17258 3782
rect 16950 3771 17258 3780
rect 21950 3836 22258 3845
rect 21950 3834 21956 3836
rect 22012 3834 22036 3836
rect 22092 3834 22116 3836
rect 22172 3834 22196 3836
rect 22252 3834 22258 3836
rect 22012 3782 22014 3834
rect 22194 3782 22196 3834
rect 21950 3780 21956 3782
rect 22012 3780 22036 3782
rect 22092 3780 22116 3782
rect 22172 3780 22196 3782
rect 22252 3780 22258 3782
rect 21950 3771 22258 3780
rect 26950 3836 27258 3845
rect 26950 3834 26956 3836
rect 27012 3834 27036 3836
rect 27092 3834 27116 3836
rect 27172 3834 27196 3836
rect 27252 3834 27258 3836
rect 27012 3782 27014 3834
rect 27194 3782 27196 3834
rect 26950 3780 26956 3782
rect 27012 3780 27036 3782
rect 27092 3780 27116 3782
rect 27172 3780 27196 3782
rect 27252 3780 27258 3782
rect 26950 3771 27258 3780
rect 31950 3836 32258 3845
rect 31950 3834 31956 3836
rect 32012 3834 32036 3836
rect 32092 3834 32116 3836
rect 32172 3834 32196 3836
rect 32252 3834 32258 3836
rect 32012 3782 32014 3834
rect 32194 3782 32196 3834
rect 31950 3780 31956 3782
rect 32012 3780 32036 3782
rect 32092 3780 32116 3782
rect 32172 3780 32196 3782
rect 32252 3780 32258 3782
rect 31950 3771 32258 3780
rect 36950 3836 37258 3845
rect 36950 3834 36956 3836
rect 37012 3834 37036 3836
rect 37092 3834 37116 3836
rect 37172 3834 37196 3836
rect 37252 3834 37258 3836
rect 37012 3782 37014 3834
rect 37194 3782 37196 3834
rect 36950 3780 36956 3782
rect 37012 3780 37036 3782
rect 37092 3780 37116 3782
rect 37172 3780 37196 3782
rect 37252 3780 37258 3782
rect 36950 3771 37258 3780
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 7610 3292 7918 3301
rect 7610 3290 7616 3292
rect 7672 3290 7696 3292
rect 7752 3290 7776 3292
rect 7832 3290 7856 3292
rect 7912 3290 7918 3292
rect 7672 3238 7674 3290
rect 7854 3238 7856 3290
rect 7610 3236 7616 3238
rect 7672 3236 7696 3238
rect 7752 3236 7776 3238
rect 7832 3236 7856 3238
rect 7912 3236 7918 3238
rect 7610 3227 7918 3236
rect 12610 3292 12918 3301
rect 12610 3290 12616 3292
rect 12672 3290 12696 3292
rect 12752 3290 12776 3292
rect 12832 3290 12856 3292
rect 12912 3290 12918 3292
rect 12672 3238 12674 3290
rect 12854 3238 12856 3290
rect 12610 3236 12616 3238
rect 12672 3236 12696 3238
rect 12752 3236 12776 3238
rect 12832 3236 12856 3238
rect 12912 3236 12918 3238
rect 12610 3227 12918 3236
rect 17610 3292 17918 3301
rect 17610 3290 17616 3292
rect 17672 3290 17696 3292
rect 17752 3290 17776 3292
rect 17832 3290 17856 3292
rect 17912 3290 17918 3292
rect 17672 3238 17674 3290
rect 17854 3238 17856 3290
rect 17610 3236 17616 3238
rect 17672 3236 17696 3238
rect 17752 3236 17776 3238
rect 17832 3236 17856 3238
rect 17912 3236 17918 3238
rect 17610 3227 17918 3236
rect 22610 3292 22918 3301
rect 22610 3290 22616 3292
rect 22672 3290 22696 3292
rect 22752 3290 22776 3292
rect 22832 3290 22856 3292
rect 22912 3290 22918 3292
rect 22672 3238 22674 3290
rect 22854 3238 22856 3290
rect 22610 3236 22616 3238
rect 22672 3236 22696 3238
rect 22752 3236 22776 3238
rect 22832 3236 22856 3238
rect 22912 3236 22918 3238
rect 22610 3227 22918 3236
rect 27610 3292 27918 3301
rect 27610 3290 27616 3292
rect 27672 3290 27696 3292
rect 27752 3290 27776 3292
rect 27832 3290 27856 3292
rect 27912 3290 27918 3292
rect 27672 3238 27674 3290
rect 27854 3238 27856 3290
rect 27610 3236 27616 3238
rect 27672 3236 27696 3238
rect 27752 3236 27776 3238
rect 27832 3236 27856 3238
rect 27912 3236 27918 3238
rect 27610 3227 27918 3236
rect 32610 3292 32918 3301
rect 32610 3290 32616 3292
rect 32672 3290 32696 3292
rect 32752 3290 32776 3292
rect 32832 3290 32856 3292
rect 32912 3290 32918 3292
rect 32672 3238 32674 3290
rect 32854 3238 32856 3290
rect 32610 3236 32616 3238
rect 32672 3236 32696 3238
rect 32752 3236 32776 3238
rect 32832 3236 32856 3238
rect 32912 3236 32918 3238
rect 32610 3227 32918 3236
rect 37610 3292 37918 3301
rect 37610 3290 37616 3292
rect 37672 3290 37696 3292
rect 37752 3290 37776 3292
rect 37832 3290 37856 3292
rect 37912 3290 37918 3292
rect 37672 3238 37674 3290
rect 37854 3238 37856 3290
rect 37610 3236 37616 3238
rect 37672 3236 37696 3238
rect 37752 3236 37776 3238
rect 37832 3236 37856 3238
rect 37912 3236 37918 3238
rect 37610 3227 37918 3236
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 6950 2748 7258 2757
rect 6950 2746 6956 2748
rect 7012 2746 7036 2748
rect 7092 2746 7116 2748
rect 7172 2746 7196 2748
rect 7252 2746 7258 2748
rect 7012 2694 7014 2746
rect 7194 2694 7196 2746
rect 6950 2692 6956 2694
rect 7012 2692 7036 2694
rect 7092 2692 7116 2694
rect 7172 2692 7196 2694
rect 7252 2692 7258 2694
rect 6950 2683 7258 2692
rect 11950 2748 12258 2757
rect 11950 2746 11956 2748
rect 12012 2746 12036 2748
rect 12092 2746 12116 2748
rect 12172 2746 12196 2748
rect 12252 2746 12258 2748
rect 12012 2694 12014 2746
rect 12194 2694 12196 2746
rect 11950 2692 11956 2694
rect 12012 2692 12036 2694
rect 12092 2692 12116 2694
rect 12172 2692 12196 2694
rect 12252 2692 12258 2694
rect 11950 2683 12258 2692
rect 16950 2748 17258 2757
rect 16950 2746 16956 2748
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17252 2746 17258 2748
rect 17012 2694 17014 2746
rect 17194 2694 17196 2746
rect 16950 2692 16956 2694
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 17252 2692 17258 2694
rect 16950 2683 17258 2692
rect 21950 2748 22258 2757
rect 21950 2746 21956 2748
rect 22012 2746 22036 2748
rect 22092 2746 22116 2748
rect 22172 2746 22196 2748
rect 22252 2746 22258 2748
rect 22012 2694 22014 2746
rect 22194 2694 22196 2746
rect 21950 2692 21956 2694
rect 22012 2692 22036 2694
rect 22092 2692 22116 2694
rect 22172 2692 22196 2694
rect 22252 2692 22258 2694
rect 21950 2683 22258 2692
rect 26950 2748 27258 2757
rect 26950 2746 26956 2748
rect 27012 2746 27036 2748
rect 27092 2746 27116 2748
rect 27172 2746 27196 2748
rect 27252 2746 27258 2748
rect 27012 2694 27014 2746
rect 27194 2694 27196 2746
rect 26950 2692 26956 2694
rect 27012 2692 27036 2694
rect 27092 2692 27116 2694
rect 27172 2692 27196 2694
rect 27252 2692 27258 2694
rect 26950 2683 27258 2692
rect 31950 2748 32258 2757
rect 31950 2746 31956 2748
rect 32012 2746 32036 2748
rect 32092 2746 32116 2748
rect 32172 2746 32196 2748
rect 32252 2746 32258 2748
rect 32012 2694 32014 2746
rect 32194 2694 32196 2746
rect 31950 2692 31956 2694
rect 32012 2692 32036 2694
rect 32092 2692 32116 2694
rect 32172 2692 32196 2694
rect 32252 2692 32258 2694
rect 31950 2683 32258 2692
rect 36950 2748 37258 2757
rect 36950 2746 36956 2748
rect 37012 2746 37036 2748
rect 37092 2746 37116 2748
rect 37172 2746 37196 2748
rect 37252 2746 37258 2748
rect 37012 2694 37014 2746
rect 37194 2694 37196 2746
rect 36950 2692 36956 2694
rect 37012 2692 37036 2694
rect 37092 2692 37116 2694
rect 37172 2692 37196 2694
rect 37252 2692 37258 2694
rect 36950 2683 37258 2692
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 7610 2204 7918 2213
rect 7610 2202 7616 2204
rect 7672 2202 7696 2204
rect 7752 2202 7776 2204
rect 7832 2202 7856 2204
rect 7912 2202 7918 2204
rect 7672 2150 7674 2202
rect 7854 2150 7856 2202
rect 7610 2148 7616 2150
rect 7672 2148 7696 2150
rect 7752 2148 7776 2150
rect 7832 2148 7856 2150
rect 7912 2148 7918 2150
rect 7610 2139 7918 2148
rect 12610 2204 12918 2213
rect 12610 2202 12616 2204
rect 12672 2202 12696 2204
rect 12752 2202 12776 2204
rect 12832 2202 12856 2204
rect 12912 2202 12918 2204
rect 12672 2150 12674 2202
rect 12854 2150 12856 2202
rect 12610 2148 12616 2150
rect 12672 2148 12696 2150
rect 12752 2148 12776 2150
rect 12832 2148 12856 2150
rect 12912 2148 12918 2150
rect 12610 2139 12918 2148
rect 17610 2204 17918 2213
rect 17610 2202 17616 2204
rect 17672 2202 17696 2204
rect 17752 2202 17776 2204
rect 17832 2202 17856 2204
rect 17912 2202 17918 2204
rect 17672 2150 17674 2202
rect 17854 2150 17856 2202
rect 17610 2148 17616 2150
rect 17672 2148 17696 2150
rect 17752 2148 17776 2150
rect 17832 2148 17856 2150
rect 17912 2148 17918 2150
rect 17610 2139 17918 2148
rect 22610 2204 22918 2213
rect 22610 2202 22616 2204
rect 22672 2202 22696 2204
rect 22752 2202 22776 2204
rect 22832 2202 22856 2204
rect 22912 2202 22918 2204
rect 22672 2150 22674 2202
rect 22854 2150 22856 2202
rect 22610 2148 22616 2150
rect 22672 2148 22696 2150
rect 22752 2148 22776 2150
rect 22832 2148 22856 2150
rect 22912 2148 22918 2150
rect 22610 2139 22918 2148
rect 27610 2204 27918 2213
rect 27610 2202 27616 2204
rect 27672 2202 27696 2204
rect 27752 2202 27776 2204
rect 27832 2202 27856 2204
rect 27912 2202 27918 2204
rect 27672 2150 27674 2202
rect 27854 2150 27856 2202
rect 27610 2148 27616 2150
rect 27672 2148 27696 2150
rect 27752 2148 27776 2150
rect 27832 2148 27856 2150
rect 27912 2148 27918 2150
rect 27610 2139 27918 2148
rect 32610 2204 32918 2213
rect 32610 2202 32616 2204
rect 32672 2202 32696 2204
rect 32752 2202 32776 2204
rect 32832 2202 32856 2204
rect 32912 2202 32918 2204
rect 32672 2150 32674 2202
rect 32854 2150 32856 2202
rect 32610 2148 32616 2150
rect 32672 2148 32696 2150
rect 32752 2148 32776 2150
rect 32832 2148 32856 2150
rect 32912 2148 32918 2150
rect 32610 2139 32918 2148
rect 37610 2204 37918 2213
rect 37610 2202 37616 2204
rect 37672 2202 37696 2204
rect 37752 2202 37776 2204
rect 37832 2202 37856 2204
rect 37912 2202 37918 2204
rect 37672 2150 37674 2202
rect 37854 2150 37856 2202
rect 37610 2148 37616 2150
rect 37672 2148 37696 2150
rect 37752 2148 37776 2150
rect 37832 2148 37856 2150
rect 37912 2148 37918 2150
rect 37610 2139 37918 2148
<< via2 >>
rect 1956 37562 2012 37564
rect 2036 37562 2092 37564
rect 2116 37562 2172 37564
rect 2196 37562 2252 37564
rect 1956 37510 2002 37562
rect 2002 37510 2012 37562
rect 2036 37510 2066 37562
rect 2066 37510 2078 37562
rect 2078 37510 2092 37562
rect 2116 37510 2130 37562
rect 2130 37510 2142 37562
rect 2142 37510 2172 37562
rect 2196 37510 2206 37562
rect 2206 37510 2252 37562
rect 1956 37508 2012 37510
rect 2036 37508 2092 37510
rect 2116 37508 2172 37510
rect 2196 37508 2252 37510
rect 6956 37562 7012 37564
rect 7036 37562 7092 37564
rect 7116 37562 7172 37564
rect 7196 37562 7252 37564
rect 6956 37510 7002 37562
rect 7002 37510 7012 37562
rect 7036 37510 7066 37562
rect 7066 37510 7078 37562
rect 7078 37510 7092 37562
rect 7116 37510 7130 37562
rect 7130 37510 7142 37562
rect 7142 37510 7172 37562
rect 7196 37510 7206 37562
rect 7206 37510 7252 37562
rect 6956 37508 7012 37510
rect 7036 37508 7092 37510
rect 7116 37508 7172 37510
rect 7196 37508 7252 37510
rect 11956 37562 12012 37564
rect 12036 37562 12092 37564
rect 12116 37562 12172 37564
rect 12196 37562 12252 37564
rect 11956 37510 12002 37562
rect 12002 37510 12012 37562
rect 12036 37510 12066 37562
rect 12066 37510 12078 37562
rect 12078 37510 12092 37562
rect 12116 37510 12130 37562
rect 12130 37510 12142 37562
rect 12142 37510 12172 37562
rect 12196 37510 12206 37562
rect 12206 37510 12252 37562
rect 11956 37508 12012 37510
rect 12036 37508 12092 37510
rect 12116 37508 12172 37510
rect 12196 37508 12252 37510
rect 16956 37562 17012 37564
rect 17036 37562 17092 37564
rect 17116 37562 17172 37564
rect 17196 37562 17252 37564
rect 16956 37510 17002 37562
rect 17002 37510 17012 37562
rect 17036 37510 17066 37562
rect 17066 37510 17078 37562
rect 17078 37510 17092 37562
rect 17116 37510 17130 37562
rect 17130 37510 17142 37562
rect 17142 37510 17172 37562
rect 17196 37510 17206 37562
rect 17206 37510 17252 37562
rect 16956 37508 17012 37510
rect 17036 37508 17092 37510
rect 17116 37508 17172 37510
rect 17196 37508 17252 37510
rect 21956 37562 22012 37564
rect 22036 37562 22092 37564
rect 22116 37562 22172 37564
rect 22196 37562 22252 37564
rect 21956 37510 22002 37562
rect 22002 37510 22012 37562
rect 22036 37510 22066 37562
rect 22066 37510 22078 37562
rect 22078 37510 22092 37562
rect 22116 37510 22130 37562
rect 22130 37510 22142 37562
rect 22142 37510 22172 37562
rect 22196 37510 22206 37562
rect 22206 37510 22252 37562
rect 21956 37508 22012 37510
rect 22036 37508 22092 37510
rect 22116 37508 22172 37510
rect 22196 37508 22252 37510
rect 26956 37562 27012 37564
rect 27036 37562 27092 37564
rect 27116 37562 27172 37564
rect 27196 37562 27252 37564
rect 26956 37510 27002 37562
rect 27002 37510 27012 37562
rect 27036 37510 27066 37562
rect 27066 37510 27078 37562
rect 27078 37510 27092 37562
rect 27116 37510 27130 37562
rect 27130 37510 27142 37562
rect 27142 37510 27172 37562
rect 27196 37510 27206 37562
rect 27206 37510 27252 37562
rect 26956 37508 27012 37510
rect 27036 37508 27092 37510
rect 27116 37508 27172 37510
rect 27196 37508 27252 37510
rect 31956 37562 32012 37564
rect 32036 37562 32092 37564
rect 32116 37562 32172 37564
rect 32196 37562 32252 37564
rect 31956 37510 32002 37562
rect 32002 37510 32012 37562
rect 32036 37510 32066 37562
rect 32066 37510 32078 37562
rect 32078 37510 32092 37562
rect 32116 37510 32130 37562
rect 32130 37510 32142 37562
rect 32142 37510 32172 37562
rect 32196 37510 32206 37562
rect 32206 37510 32252 37562
rect 31956 37508 32012 37510
rect 32036 37508 32092 37510
rect 32116 37508 32172 37510
rect 32196 37508 32252 37510
rect 36956 37562 37012 37564
rect 37036 37562 37092 37564
rect 37116 37562 37172 37564
rect 37196 37562 37252 37564
rect 36956 37510 37002 37562
rect 37002 37510 37012 37562
rect 37036 37510 37066 37562
rect 37066 37510 37078 37562
rect 37078 37510 37092 37562
rect 37116 37510 37130 37562
rect 37130 37510 37142 37562
rect 37142 37510 37172 37562
rect 37196 37510 37206 37562
rect 37206 37510 37252 37562
rect 36956 37508 37012 37510
rect 37036 37508 37092 37510
rect 37116 37508 37172 37510
rect 37196 37508 37252 37510
rect 2616 37018 2672 37020
rect 2696 37018 2752 37020
rect 2776 37018 2832 37020
rect 2856 37018 2912 37020
rect 2616 36966 2662 37018
rect 2662 36966 2672 37018
rect 2696 36966 2726 37018
rect 2726 36966 2738 37018
rect 2738 36966 2752 37018
rect 2776 36966 2790 37018
rect 2790 36966 2802 37018
rect 2802 36966 2832 37018
rect 2856 36966 2866 37018
rect 2866 36966 2912 37018
rect 2616 36964 2672 36966
rect 2696 36964 2752 36966
rect 2776 36964 2832 36966
rect 2856 36964 2912 36966
rect 7616 37018 7672 37020
rect 7696 37018 7752 37020
rect 7776 37018 7832 37020
rect 7856 37018 7912 37020
rect 7616 36966 7662 37018
rect 7662 36966 7672 37018
rect 7696 36966 7726 37018
rect 7726 36966 7738 37018
rect 7738 36966 7752 37018
rect 7776 36966 7790 37018
rect 7790 36966 7802 37018
rect 7802 36966 7832 37018
rect 7856 36966 7866 37018
rect 7866 36966 7912 37018
rect 7616 36964 7672 36966
rect 7696 36964 7752 36966
rect 7776 36964 7832 36966
rect 7856 36964 7912 36966
rect 12616 37018 12672 37020
rect 12696 37018 12752 37020
rect 12776 37018 12832 37020
rect 12856 37018 12912 37020
rect 12616 36966 12662 37018
rect 12662 36966 12672 37018
rect 12696 36966 12726 37018
rect 12726 36966 12738 37018
rect 12738 36966 12752 37018
rect 12776 36966 12790 37018
rect 12790 36966 12802 37018
rect 12802 36966 12832 37018
rect 12856 36966 12866 37018
rect 12866 36966 12912 37018
rect 12616 36964 12672 36966
rect 12696 36964 12752 36966
rect 12776 36964 12832 36966
rect 12856 36964 12912 36966
rect 17616 37018 17672 37020
rect 17696 37018 17752 37020
rect 17776 37018 17832 37020
rect 17856 37018 17912 37020
rect 17616 36966 17662 37018
rect 17662 36966 17672 37018
rect 17696 36966 17726 37018
rect 17726 36966 17738 37018
rect 17738 36966 17752 37018
rect 17776 36966 17790 37018
rect 17790 36966 17802 37018
rect 17802 36966 17832 37018
rect 17856 36966 17866 37018
rect 17866 36966 17912 37018
rect 17616 36964 17672 36966
rect 17696 36964 17752 36966
rect 17776 36964 17832 36966
rect 17856 36964 17912 36966
rect 22616 37018 22672 37020
rect 22696 37018 22752 37020
rect 22776 37018 22832 37020
rect 22856 37018 22912 37020
rect 22616 36966 22662 37018
rect 22662 36966 22672 37018
rect 22696 36966 22726 37018
rect 22726 36966 22738 37018
rect 22738 36966 22752 37018
rect 22776 36966 22790 37018
rect 22790 36966 22802 37018
rect 22802 36966 22832 37018
rect 22856 36966 22866 37018
rect 22866 36966 22912 37018
rect 22616 36964 22672 36966
rect 22696 36964 22752 36966
rect 22776 36964 22832 36966
rect 22856 36964 22912 36966
rect 27616 37018 27672 37020
rect 27696 37018 27752 37020
rect 27776 37018 27832 37020
rect 27856 37018 27912 37020
rect 27616 36966 27662 37018
rect 27662 36966 27672 37018
rect 27696 36966 27726 37018
rect 27726 36966 27738 37018
rect 27738 36966 27752 37018
rect 27776 36966 27790 37018
rect 27790 36966 27802 37018
rect 27802 36966 27832 37018
rect 27856 36966 27866 37018
rect 27866 36966 27912 37018
rect 27616 36964 27672 36966
rect 27696 36964 27752 36966
rect 27776 36964 27832 36966
rect 27856 36964 27912 36966
rect 32616 37018 32672 37020
rect 32696 37018 32752 37020
rect 32776 37018 32832 37020
rect 32856 37018 32912 37020
rect 32616 36966 32662 37018
rect 32662 36966 32672 37018
rect 32696 36966 32726 37018
rect 32726 36966 32738 37018
rect 32738 36966 32752 37018
rect 32776 36966 32790 37018
rect 32790 36966 32802 37018
rect 32802 36966 32832 37018
rect 32856 36966 32866 37018
rect 32866 36966 32912 37018
rect 32616 36964 32672 36966
rect 32696 36964 32752 36966
rect 32776 36964 32832 36966
rect 32856 36964 32912 36966
rect 37616 37018 37672 37020
rect 37696 37018 37752 37020
rect 37776 37018 37832 37020
rect 37856 37018 37912 37020
rect 37616 36966 37662 37018
rect 37662 36966 37672 37018
rect 37696 36966 37726 37018
rect 37726 36966 37738 37018
rect 37738 36966 37752 37018
rect 37776 36966 37790 37018
rect 37790 36966 37802 37018
rect 37802 36966 37832 37018
rect 37856 36966 37866 37018
rect 37866 36966 37912 37018
rect 37616 36964 37672 36966
rect 37696 36964 37752 36966
rect 37776 36964 37832 36966
rect 37856 36964 37912 36966
rect 1956 36474 2012 36476
rect 2036 36474 2092 36476
rect 2116 36474 2172 36476
rect 2196 36474 2252 36476
rect 1956 36422 2002 36474
rect 2002 36422 2012 36474
rect 2036 36422 2066 36474
rect 2066 36422 2078 36474
rect 2078 36422 2092 36474
rect 2116 36422 2130 36474
rect 2130 36422 2142 36474
rect 2142 36422 2172 36474
rect 2196 36422 2206 36474
rect 2206 36422 2252 36474
rect 1956 36420 2012 36422
rect 2036 36420 2092 36422
rect 2116 36420 2172 36422
rect 2196 36420 2252 36422
rect 6956 36474 7012 36476
rect 7036 36474 7092 36476
rect 7116 36474 7172 36476
rect 7196 36474 7252 36476
rect 6956 36422 7002 36474
rect 7002 36422 7012 36474
rect 7036 36422 7066 36474
rect 7066 36422 7078 36474
rect 7078 36422 7092 36474
rect 7116 36422 7130 36474
rect 7130 36422 7142 36474
rect 7142 36422 7172 36474
rect 7196 36422 7206 36474
rect 7206 36422 7252 36474
rect 6956 36420 7012 36422
rect 7036 36420 7092 36422
rect 7116 36420 7172 36422
rect 7196 36420 7252 36422
rect 11956 36474 12012 36476
rect 12036 36474 12092 36476
rect 12116 36474 12172 36476
rect 12196 36474 12252 36476
rect 11956 36422 12002 36474
rect 12002 36422 12012 36474
rect 12036 36422 12066 36474
rect 12066 36422 12078 36474
rect 12078 36422 12092 36474
rect 12116 36422 12130 36474
rect 12130 36422 12142 36474
rect 12142 36422 12172 36474
rect 12196 36422 12206 36474
rect 12206 36422 12252 36474
rect 11956 36420 12012 36422
rect 12036 36420 12092 36422
rect 12116 36420 12172 36422
rect 12196 36420 12252 36422
rect 16956 36474 17012 36476
rect 17036 36474 17092 36476
rect 17116 36474 17172 36476
rect 17196 36474 17252 36476
rect 16956 36422 17002 36474
rect 17002 36422 17012 36474
rect 17036 36422 17066 36474
rect 17066 36422 17078 36474
rect 17078 36422 17092 36474
rect 17116 36422 17130 36474
rect 17130 36422 17142 36474
rect 17142 36422 17172 36474
rect 17196 36422 17206 36474
rect 17206 36422 17252 36474
rect 16956 36420 17012 36422
rect 17036 36420 17092 36422
rect 17116 36420 17172 36422
rect 17196 36420 17252 36422
rect 21956 36474 22012 36476
rect 22036 36474 22092 36476
rect 22116 36474 22172 36476
rect 22196 36474 22252 36476
rect 21956 36422 22002 36474
rect 22002 36422 22012 36474
rect 22036 36422 22066 36474
rect 22066 36422 22078 36474
rect 22078 36422 22092 36474
rect 22116 36422 22130 36474
rect 22130 36422 22142 36474
rect 22142 36422 22172 36474
rect 22196 36422 22206 36474
rect 22206 36422 22252 36474
rect 21956 36420 22012 36422
rect 22036 36420 22092 36422
rect 22116 36420 22172 36422
rect 22196 36420 22252 36422
rect 26956 36474 27012 36476
rect 27036 36474 27092 36476
rect 27116 36474 27172 36476
rect 27196 36474 27252 36476
rect 26956 36422 27002 36474
rect 27002 36422 27012 36474
rect 27036 36422 27066 36474
rect 27066 36422 27078 36474
rect 27078 36422 27092 36474
rect 27116 36422 27130 36474
rect 27130 36422 27142 36474
rect 27142 36422 27172 36474
rect 27196 36422 27206 36474
rect 27206 36422 27252 36474
rect 26956 36420 27012 36422
rect 27036 36420 27092 36422
rect 27116 36420 27172 36422
rect 27196 36420 27252 36422
rect 31956 36474 32012 36476
rect 32036 36474 32092 36476
rect 32116 36474 32172 36476
rect 32196 36474 32252 36476
rect 31956 36422 32002 36474
rect 32002 36422 32012 36474
rect 32036 36422 32066 36474
rect 32066 36422 32078 36474
rect 32078 36422 32092 36474
rect 32116 36422 32130 36474
rect 32130 36422 32142 36474
rect 32142 36422 32172 36474
rect 32196 36422 32206 36474
rect 32206 36422 32252 36474
rect 31956 36420 32012 36422
rect 32036 36420 32092 36422
rect 32116 36420 32172 36422
rect 32196 36420 32252 36422
rect 36956 36474 37012 36476
rect 37036 36474 37092 36476
rect 37116 36474 37172 36476
rect 37196 36474 37252 36476
rect 36956 36422 37002 36474
rect 37002 36422 37012 36474
rect 37036 36422 37066 36474
rect 37066 36422 37078 36474
rect 37078 36422 37092 36474
rect 37116 36422 37130 36474
rect 37130 36422 37142 36474
rect 37142 36422 37172 36474
rect 37196 36422 37206 36474
rect 37206 36422 37252 36474
rect 36956 36420 37012 36422
rect 37036 36420 37092 36422
rect 37116 36420 37172 36422
rect 37196 36420 37252 36422
rect 2616 35930 2672 35932
rect 2696 35930 2752 35932
rect 2776 35930 2832 35932
rect 2856 35930 2912 35932
rect 2616 35878 2662 35930
rect 2662 35878 2672 35930
rect 2696 35878 2726 35930
rect 2726 35878 2738 35930
rect 2738 35878 2752 35930
rect 2776 35878 2790 35930
rect 2790 35878 2802 35930
rect 2802 35878 2832 35930
rect 2856 35878 2866 35930
rect 2866 35878 2912 35930
rect 2616 35876 2672 35878
rect 2696 35876 2752 35878
rect 2776 35876 2832 35878
rect 2856 35876 2912 35878
rect 7616 35930 7672 35932
rect 7696 35930 7752 35932
rect 7776 35930 7832 35932
rect 7856 35930 7912 35932
rect 7616 35878 7662 35930
rect 7662 35878 7672 35930
rect 7696 35878 7726 35930
rect 7726 35878 7738 35930
rect 7738 35878 7752 35930
rect 7776 35878 7790 35930
rect 7790 35878 7802 35930
rect 7802 35878 7832 35930
rect 7856 35878 7866 35930
rect 7866 35878 7912 35930
rect 7616 35876 7672 35878
rect 7696 35876 7752 35878
rect 7776 35876 7832 35878
rect 7856 35876 7912 35878
rect 12616 35930 12672 35932
rect 12696 35930 12752 35932
rect 12776 35930 12832 35932
rect 12856 35930 12912 35932
rect 12616 35878 12662 35930
rect 12662 35878 12672 35930
rect 12696 35878 12726 35930
rect 12726 35878 12738 35930
rect 12738 35878 12752 35930
rect 12776 35878 12790 35930
rect 12790 35878 12802 35930
rect 12802 35878 12832 35930
rect 12856 35878 12866 35930
rect 12866 35878 12912 35930
rect 12616 35876 12672 35878
rect 12696 35876 12752 35878
rect 12776 35876 12832 35878
rect 12856 35876 12912 35878
rect 17616 35930 17672 35932
rect 17696 35930 17752 35932
rect 17776 35930 17832 35932
rect 17856 35930 17912 35932
rect 17616 35878 17662 35930
rect 17662 35878 17672 35930
rect 17696 35878 17726 35930
rect 17726 35878 17738 35930
rect 17738 35878 17752 35930
rect 17776 35878 17790 35930
rect 17790 35878 17802 35930
rect 17802 35878 17832 35930
rect 17856 35878 17866 35930
rect 17866 35878 17912 35930
rect 17616 35876 17672 35878
rect 17696 35876 17752 35878
rect 17776 35876 17832 35878
rect 17856 35876 17912 35878
rect 22616 35930 22672 35932
rect 22696 35930 22752 35932
rect 22776 35930 22832 35932
rect 22856 35930 22912 35932
rect 22616 35878 22662 35930
rect 22662 35878 22672 35930
rect 22696 35878 22726 35930
rect 22726 35878 22738 35930
rect 22738 35878 22752 35930
rect 22776 35878 22790 35930
rect 22790 35878 22802 35930
rect 22802 35878 22832 35930
rect 22856 35878 22866 35930
rect 22866 35878 22912 35930
rect 22616 35876 22672 35878
rect 22696 35876 22752 35878
rect 22776 35876 22832 35878
rect 22856 35876 22912 35878
rect 27616 35930 27672 35932
rect 27696 35930 27752 35932
rect 27776 35930 27832 35932
rect 27856 35930 27912 35932
rect 27616 35878 27662 35930
rect 27662 35878 27672 35930
rect 27696 35878 27726 35930
rect 27726 35878 27738 35930
rect 27738 35878 27752 35930
rect 27776 35878 27790 35930
rect 27790 35878 27802 35930
rect 27802 35878 27832 35930
rect 27856 35878 27866 35930
rect 27866 35878 27912 35930
rect 27616 35876 27672 35878
rect 27696 35876 27752 35878
rect 27776 35876 27832 35878
rect 27856 35876 27912 35878
rect 32616 35930 32672 35932
rect 32696 35930 32752 35932
rect 32776 35930 32832 35932
rect 32856 35930 32912 35932
rect 32616 35878 32662 35930
rect 32662 35878 32672 35930
rect 32696 35878 32726 35930
rect 32726 35878 32738 35930
rect 32738 35878 32752 35930
rect 32776 35878 32790 35930
rect 32790 35878 32802 35930
rect 32802 35878 32832 35930
rect 32856 35878 32866 35930
rect 32866 35878 32912 35930
rect 32616 35876 32672 35878
rect 32696 35876 32752 35878
rect 32776 35876 32832 35878
rect 32856 35876 32912 35878
rect 37616 35930 37672 35932
rect 37696 35930 37752 35932
rect 37776 35930 37832 35932
rect 37856 35930 37912 35932
rect 37616 35878 37662 35930
rect 37662 35878 37672 35930
rect 37696 35878 37726 35930
rect 37726 35878 37738 35930
rect 37738 35878 37752 35930
rect 37776 35878 37790 35930
rect 37790 35878 37802 35930
rect 37802 35878 37832 35930
rect 37856 35878 37866 35930
rect 37866 35878 37912 35930
rect 37616 35876 37672 35878
rect 37696 35876 37752 35878
rect 37776 35876 37832 35878
rect 37856 35876 37912 35878
rect 1956 35386 2012 35388
rect 2036 35386 2092 35388
rect 2116 35386 2172 35388
rect 2196 35386 2252 35388
rect 1956 35334 2002 35386
rect 2002 35334 2012 35386
rect 2036 35334 2066 35386
rect 2066 35334 2078 35386
rect 2078 35334 2092 35386
rect 2116 35334 2130 35386
rect 2130 35334 2142 35386
rect 2142 35334 2172 35386
rect 2196 35334 2206 35386
rect 2206 35334 2252 35386
rect 1956 35332 2012 35334
rect 2036 35332 2092 35334
rect 2116 35332 2172 35334
rect 2196 35332 2252 35334
rect 6956 35386 7012 35388
rect 7036 35386 7092 35388
rect 7116 35386 7172 35388
rect 7196 35386 7252 35388
rect 6956 35334 7002 35386
rect 7002 35334 7012 35386
rect 7036 35334 7066 35386
rect 7066 35334 7078 35386
rect 7078 35334 7092 35386
rect 7116 35334 7130 35386
rect 7130 35334 7142 35386
rect 7142 35334 7172 35386
rect 7196 35334 7206 35386
rect 7206 35334 7252 35386
rect 6956 35332 7012 35334
rect 7036 35332 7092 35334
rect 7116 35332 7172 35334
rect 7196 35332 7252 35334
rect 11956 35386 12012 35388
rect 12036 35386 12092 35388
rect 12116 35386 12172 35388
rect 12196 35386 12252 35388
rect 11956 35334 12002 35386
rect 12002 35334 12012 35386
rect 12036 35334 12066 35386
rect 12066 35334 12078 35386
rect 12078 35334 12092 35386
rect 12116 35334 12130 35386
rect 12130 35334 12142 35386
rect 12142 35334 12172 35386
rect 12196 35334 12206 35386
rect 12206 35334 12252 35386
rect 11956 35332 12012 35334
rect 12036 35332 12092 35334
rect 12116 35332 12172 35334
rect 12196 35332 12252 35334
rect 16956 35386 17012 35388
rect 17036 35386 17092 35388
rect 17116 35386 17172 35388
rect 17196 35386 17252 35388
rect 16956 35334 17002 35386
rect 17002 35334 17012 35386
rect 17036 35334 17066 35386
rect 17066 35334 17078 35386
rect 17078 35334 17092 35386
rect 17116 35334 17130 35386
rect 17130 35334 17142 35386
rect 17142 35334 17172 35386
rect 17196 35334 17206 35386
rect 17206 35334 17252 35386
rect 16956 35332 17012 35334
rect 17036 35332 17092 35334
rect 17116 35332 17172 35334
rect 17196 35332 17252 35334
rect 21956 35386 22012 35388
rect 22036 35386 22092 35388
rect 22116 35386 22172 35388
rect 22196 35386 22252 35388
rect 21956 35334 22002 35386
rect 22002 35334 22012 35386
rect 22036 35334 22066 35386
rect 22066 35334 22078 35386
rect 22078 35334 22092 35386
rect 22116 35334 22130 35386
rect 22130 35334 22142 35386
rect 22142 35334 22172 35386
rect 22196 35334 22206 35386
rect 22206 35334 22252 35386
rect 21956 35332 22012 35334
rect 22036 35332 22092 35334
rect 22116 35332 22172 35334
rect 22196 35332 22252 35334
rect 26956 35386 27012 35388
rect 27036 35386 27092 35388
rect 27116 35386 27172 35388
rect 27196 35386 27252 35388
rect 26956 35334 27002 35386
rect 27002 35334 27012 35386
rect 27036 35334 27066 35386
rect 27066 35334 27078 35386
rect 27078 35334 27092 35386
rect 27116 35334 27130 35386
rect 27130 35334 27142 35386
rect 27142 35334 27172 35386
rect 27196 35334 27206 35386
rect 27206 35334 27252 35386
rect 26956 35332 27012 35334
rect 27036 35332 27092 35334
rect 27116 35332 27172 35334
rect 27196 35332 27252 35334
rect 31956 35386 32012 35388
rect 32036 35386 32092 35388
rect 32116 35386 32172 35388
rect 32196 35386 32252 35388
rect 31956 35334 32002 35386
rect 32002 35334 32012 35386
rect 32036 35334 32066 35386
rect 32066 35334 32078 35386
rect 32078 35334 32092 35386
rect 32116 35334 32130 35386
rect 32130 35334 32142 35386
rect 32142 35334 32172 35386
rect 32196 35334 32206 35386
rect 32206 35334 32252 35386
rect 31956 35332 32012 35334
rect 32036 35332 32092 35334
rect 32116 35332 32172 35334
rect 32196 35332 32252 35334
rect 36956 35386 37012 35388
rect 37036 35386 37092 35388
rect 37116 35386 37172 35388
rect 37196 35386 37252 35388
rect 36956 35334 37002 35386
rect 37002 35334 37012 35386
rect 37036 35334 37066 35386
rect 37066 35334 37078 35386
rect 37078 35334 37092 35386
rect 37116 35334 37130 35386
rect 37130 35334 37142 35386
rect 37142 35334 37172 35386
rect 37196 35334 37206 35386
rect 37206 35334 37252 35386
rect 36956 35332 37012 35334
rect 37036 35332 37092 35334
rect 37116 35332 37172 35334
rect 37196 35332 37252 35334
rect 2616 34842 2672 34844
rect 2696 34842 2752 34844
rect 2776 34842 2832 34844
rect 2856 34842 2912 34844
rect 2616 34790 2662 34842
rect 2662 34790 2672 34842
rect 2696 34790 2726 34842
rect 2726 34790 2738 34842
rect 2738 34790 2752 34842
rect 2776 34790 2790 34842
rect 2790 34790 2802 34842
rect 2802 34790 2832 34842
rect 2856 34790 2866 34842
rect 2866 34790 2912 34842
rect 2616 34788 2672 34790
rect 2696 34788 2752 34790
rect 2776 34788 2832 34790
rect 2856 34788 2912 34790
rect 7616 34842 7672 34844
rect 7696 34842 7752 34844
rect 7776 34842 7832 34844
rect 7856 34842 7912 34844
rect 7616 34790 7662 34842
rect 7662 34790 7672 34842
rect 7696 34790 7726 34842
rect 7726 34790 7738 34842
rect 7738 34790 7752 34842
rect 7776 34790 7790 34842
rect 7790 34790 7802 34842
rect 7802 34790 7832 34842
rect 7856 34790 7866 34842
rect 7866 34790 7912 34842
rect 7616 34788 7672 34790
rect 7696 34788 7752 34790
rect 7776 34788 7832 34790
rect 7856 34788 7912 34790
rect 12616 34842 12672 34844
rect 12696 34842 12752 34844
rect 12776 34842 12832 34844
rect 12856 34842 12912 34844
rect 12616 34790 12662 34842
rect 12662 34790 12672 34842
rect 12696 34790 12726 34842
rect 12726 34790 12738 34842
rect 12738 34790 12752 34842
rect 12776 34790 12790 34842
rect 12790 34790 12802 34842
rect 12802 34790 12832 34842
rect 12856 34790 12866 34842
rect 12866 34790 12912 34842
rect 12616 34788 12672 34790
rect 12696 34788 12752 34790
rect 12776 34788 12832 34790
rect 12856 34788 12912 34790
rect 17616 34842 17672 34844
rect 17696 34842 17752 34844
rect 17776 34842 17832 34844
rect 17856 34842 17912 34844
rect 17616 34790 17662 34842
rect 17662 34790 17672 34842
rect 17696 34790 17726 34842
rect 17726 34790 17738 34842
rect 17738 34790 17752 34842
rect 17776 34790 17790 34842
rect 17790 34790 17802 34842
rect 17802 34790 17832 34842
rect 17856 34790 17866 34842
rect 17866 34790 17912 34842
rect 17616 34788 17672 34790
rect 17696 34788 17752 34790
rect 17776 34788 17832 34790
rect 17856 34788 17912 34790
rect 22616 34842 22672 34844
rect 22696 34842 22752 34844
rect 22776 34842 22832 34844
rect 22856 34842 22912 34844
rect 22616 34790 22662 34842
rect 22662 34790 22672 34842
rect 22696 34790 22726 34842
rect 22726 34790 22738 34842
rect 22738 34790 22752 34842
rect 22776 34790 22790 34842
rect 22790 34790 22802 34842
rect 22802 34790 22832 34842
rect 22856 34790 22866 34842
rect 22866 34790 22912 34842
rect 22616 34788 22672 34790
rect 22696 34788 22752 34790
rect 22776 34788 22832 34790
rect 22856 34788 22912 34790
rect 27616 34842 27672 34844
rect 27696 34842 27752 34844
rect 27776 34842 27832 34844
rect 27856 34842 27912 34844
rect 27616 34790 27662 34842
rect 27662 34790 27672 34842
rect 27696 34790 27726 34842
rect 27726 34790 27738 34842
rect 27738 34790 27752 34842
rect 27776 34790 27790 34842
rect 27790 34790 27802 34842
rect 27802 34790 27832 34842
rect 27856 34790 27866 34842
rect 27866 34790 27912 34842
rect 27616 34788 27672 34790
rect 27696 34788 27752 34790
rect 27776 34788 27832 34790
rect 27856 34788 27912 34790
rect 32616 34842 32672 34844
rect 32696 34842 32752 34844
rect 32776 34842 32832 34844
rect 32856 34842 32912 34844
rect 32616 34790 32662 34842
rect 32662 34790 32672 34842
rect 32696 34790 32726 34842
rect 32726 34790 32738 34842
rect 32738 34790 32752 34842
rect 32776 34790 32790 34842
rect 32790 34790 32802 34842
rect 32802 34790 32832 34842
rect 32856 34790 32866 34842
rect 32866 34790 32912 34842
rect 32616 34788 32672 34790
rect 32696 34788 32752 34790
rect 32776 34788 32832 34790
rect 32856 34788 32912 34790
rect 37616 34842 37672 34844
rect 37696 34842 37752 34844
rect 37776 34842 37832 34844
rect 37856 34842 37912 34844
rect 37616 34790 37662 34842
rect 37662 34790 37672 34842
rect 37696 34790 37726 34842
rect 37726 34790 37738 34842
rect 37738 34790 37752 34842
rect 37776 34790 37790 34842
rect 37790 34790 37802 34842
rect 37802 34790 37832 34842
rect 37856 34790 37866 34842
rect 37866 34790 37912 34842
rect 37616 34788 37672 34790
rect 37696 34788 37752 34790
rect 37776 34788 37832 34790
rect 37856 34788 37912 34790
rect 1956 34298 2012 34300
rect 2036 34298 2092 34300
rect 2116 34298 2172 34300
rect 2196 34298 2252 34300
rect 1956 34246 2002 34298
rect 2002 34246 2012 34298
rect 2036 34246 2066 34298
rect 2066 34246 2078 34298
rect 2078 34246 2092 34298
rect 2116 34246 2130 34298
rect 2130 34246 2142 34298
rect 2142 34246 2172 34298
rect 2196 34246 2206 34298
rect 2206 34246 2252 34298
rect 1956 34244 2012 34246
rect 2036 34244 2092 34246
rect 2116 34244 2172 34246
rect 2196 34244 2252 34246
rect 6956 34298 7012 34300
rect 7036 34298 7092 34300
rect 7116 34298 7172 34300
rect 7196 34298 7252 34300
rect 6956 34246 7002 34298
rect 7002 34246 7012 34298
rect 7036 34246 7066 34298
rect 7066 34246 7078 34298
rect 7078 34246 7092 34298
rect 7116 34246 7130 34298
rect 7130 34246 7142 34298
rect 7142 34246 7172 34298
rect 7196 34246 7206 34298
rect 7206 34246 7252 34298
rect 6956 34244 7012 34246
rect 7036 34244 7092 34246
rect 7116 34244 7172 34246
rect 7196 34244 7252 34246
rect 11956 34298 12012 34300
rect 12036 34298 12092 34300
rect 12116 34298 12172 34300
rect 12196 34298 12252 34300
rect 11956 34246 12002 34298
rect 12002 34246 12012 34298
rect 12036 34246 12066 34298
rect 12066 34246 12078 34298
rect 12078 34246 12092 34298
rect 12116 34246 12130 34298
rect 12130 34246 12142 34298
rect 12142 34246 12172 34298
rect 12196 34246 12206 34298
rect 12206 34246 12252 34298
rect 11956 34244 12012 34246
rect 12036 34244 12092 34246
rect 12116 34244 12172 34246
rect 12196 34244 12252 34246
rect 16956 34298 17012 34300
rect 17036 34298 17092 34300
rect 17116 34298 17172 34300
rect 17196 34298 17252 34300
rect 16956 34246 17002 34298
rect 17002 34246 17012 34298
rect 17036 34246 17066 34298
rect 17066 34246 17078 34298
rect 17078 34246 17092 34298
rect 17116 34246 17130 34298
rect 17130 34246 17142 34298
rect 17142 34246 17172 34298
rect 17196 34246 17206 34298
rect 17206 34246 17252 34298
rect 16956 34244 17012 34246
rect 17036 34244 17092 34246
rect 17116 34244 17172 34246
rect 17196 34244 17252 34246
rect 21956 34298 22012 34300
rect 22036 34298 22092 34300
rect 22116 34298 22172 34300
rect 22196 34298 22252 34300
rect 21956 34246 22002 34298
rect 22002 34246 22012 34298
rect 22036 34246 22066 34298
rect 22066 34246 22078 34298
rect 22078 34246 22092 34298
rect 22116 34246 22130 34298
rect 22130 34246 22142 34298
rect 22142 34246 22172 34298
rect 22196 34246 22206 34298
rect 22206 34246 22252 34298
rect 21956 34244 22012 34246
rect 22036 34244 22092 34246
rect 22116 34244 22172 34246
rect 22196 34244 22252 34246
rect 26956 34298 27012 34300
rect 27036 34298 27092 34300
rect 27116 34298 27172 34300
rect 27196 34298 27252 34300
rect 26956 34246 27002 34298
rect 27002 34246 27012 34298
rect 27036 34246 27066 34298
rect 27066 34246 27078 34298
rect 27078 34246 27092 34298
rect 27116 34246 27130 34298
rect 27130 34246 27142 34298
rect 27142 34246 27172 34298
rect 27196 34246 27206 34298
rect 27206 34246 27252 34298
rect 26956 34244 27012 34246
rect 27036 34244 27092 34246
rect 27116 34244 27172 34246
rect 27196 34244 27252 34246
rect 31956 34298 32012 34300
rect 32036 34298 32092 34300
rect 32116 34298 32172 34300
rect 32196 34298 32252 34300
rect 31956 34246 32002 34298
rect 32002 34246 32012 34298
rect 32036 34246 32066 34298
rect 32066 34246 32078 34298
rect 32078 34246 32092 34298
rect 32116 34246 32130 34298
rect 32130 34246 32142 34298
rect 32142 34246 32172 34298
rect 32196 34246 32206 34298
rect 32206 34246 32252 34298
rect 31956 34244 32012 34246
rect 32036 34244 32092 34246
rect 32116 34244 32172 34246
rect 32196 34244 32252 34246
rect 36956 34298 37012 34300
rect 37036 34298 37092 34300
rect 37116 34298 37172 34300
rect 37196 34298 37252 34300
rect 36956 34246 37002 34298
rect 37002 34246 37012 34298
rect 37036 34246 37066 34298
rect 37066 34246 37078 34298
rect 37078 34246 37092 34298
rect 37116 34246 37130 34298
rect 37130 34246 37142 34298
rect 37142 34246 37172 34298
rect 37196 34246 37206 34298
rect 37206 34246 37252 34298
rect 36956 34244 37012 34246
rect 37036 34244 37092 34246
rect 37116 34244 37172 34246
rect 37196 34244 37252 34246
rect 2616 33754 2672 33756
rect 2696 33754 2752 33756
rect 2776 33754 2832 33756
rect 2856 33754 2912 33756
rect 2616 33702 2662 33754
rect 2662 33702 2672 33754
rect 2696 33702 2726 33754
rect 2726 33702 2738 33754
rect 2738 33702 2752 33754
rect 2776 33702 2790 33754
rect 2790 33702 2802 33754
rect 2802 33702 2832 33754
rect 2856 33702 2866 33754
rect 2866 33702 2912 33754
rect 2616 33700 2672 33702
rect 2696 33700 2752 33702
rect 2776 33700 2832 33702
rect 2856 33700 2912 33702
rect 7616 33754 7672 33756
rect 7696 33754 7752 33756
rect 7776 33754 7832 33756
rect 7856 33754 7912 33756
rect 7616 33702 7662 33754
rect 7662 33702 7672 33754
rect 7696 33702 7726 33754
rect 7726 33702 7738 33754
rect 7738 33702 7752 33754
rect 7776 33702 7790 33754
rect 7790 33702 7802 33754
rect 7802 33702 7832 33754
rect 7856 33702 7866 33754
rect 7866 33702 7912 33754
rect 7616 33700 7672 33702
rect 7696 33700 7752 33702
rect 7776 33700 7832 33702
rect 7856 33700 7912 33702
rect 12616 33754 12672 33756
rect 12696 33754 12752 33756
rect 12776 33754 12832 33756
rect 12856 33754 12912 33756
rect 12616 33702 12662 33754
rect 12662 33702 12672 33754
rect 12696 33702 12726 33754
rect 12726 33702 12738 33754
rect 12738 33702 12752 33754
rect 12776 33702 12790 33754
rect 12790 33702 12802 33754
rect 12802 33702 12832 33754
rect 12856 33702 12866 33754
rect 12866 33702 12912 33754
rect 12616 33700 12672 33702
rect 12696 33700 12752 33702
rect 12776 33700 12832 33702
rect 12856 33700 12912 33702
rect 17616 33754 17672 33756
rect 17696 33754 17752 33756
rect 17776 33754 17832 33756
rect 17856 33754 17912 33756
rect 17616 33702 17662 33754
rect 17662 33702 17672 33754
rect 17696 33702 17726 33754
rect 17726 33702 17738 33754
rect 17738 33702 17752 33754
rect 17776 33702 17790 33754
rect 17790 33702 17802 33754
rect 17802 33702 17832 33754
rect 17856 33702 17866 33754
rect 17866 33702 17912 33754
rect 17616 33700 17672 33702
rect 17696 33700 17752 33702
rect 17776 33700 17832 33702
rect 17856 33700 17912 33702
rect 22616 33754 22672 33756
rect 22696 33754 22752 33756
rect 22776 33754 22832 33756
rect 22856 33754 22912 33756
rect 22616 33702 22662 33754
rect 22662 33702 22672 33754
rect 22696 33702 22726 33754
rect 22726 33702 22738 33754
rect 22738 33702 22752 33754
rect 22776 33702 22790 33754
rect 22790 33702 22802 33754
rect 22802 33702 22832 33754
rect 22856 33702 22866 33754
rect 22866 33702 22912 33754
rect 22616 33700 22672 33702
rect 22696 33700 22752 33702
rect 22776 33700 22832 33702
rect 22856 33700 22912 33702
rect 27616 33754 27672 33756
rect 27696 33754 27752 33756
rect 27776 33754 27832 33756
rect 27856 33754 27912 33756
rect 27616 33702 27662 33754
rect 27662 33702 27672 33754
rect 27696 33702 27726 33754
rect 27726 33702 27738 33754
rect 27738 33702 27752 33754
rect 27776 33702 27790 33754
rect 27790 33702 27802 33754
rect 27802 33702 27832 33754
rect 27856 33702 27866 33754
rect 27866 33702 27912 33754
rect 27616 33700 27672 33702
rect 27696 33700 27752 33702
rect 27776 33700 27832 33702
rect 27856 33700 27912 33702
rect 32616 33754 32672 33756
rect 32696 33754 32752 33756
rect 32776 33754 32832 33756
rect 32856 33754 32912 33756
rect 32616 33702 32662 33754
rect 32662 33702 32672 33754
rect 32696 33702 32726 33754
rect 32726 33702 32738 33754
rect 32738 33702 32752 33754
rect 32776 33702 32790 33754
rect 32790 33702 32802 33754
rect 32802 33702 32832 33754
rect 32856 33702 32866 33754
rect 32866 33702 32912 33754
rect 32616 33700 32672 33702
rect 32696 33700 32752 33702
rect 32776 33700 32832 33702
rect 32856 33700 32912 33702
rect 37616 33754 37672 33756
rect 37696 33754 37752 33756
rect 37776 33754 37832 33756
rect 37856 33754 37912 33756
rect 37616 33702 37662 33754
rect 37662 33702 37672 33754
rect 37696 33702 37726 33754
rect 37726 33702 37738 33754
rect 37738 33702 37752 33754
rect 37776 33702 37790 33754
rect 37790 33702 37802 33754
rect 37802 33702 37832 33754
rect 37856 33702 37866 33754
rect 37866 33702 37912 33754
rect 37616 33700 37672 33702
rect 37696 33700 37752 33702
rect 37776 33700 37832 33702
rect 37856 33700 37912 33702
rect 1956 33210 2012 33212
rect 2036 33210 2092 33212
rect 2116 33210 2172 33212
rect 2196 33210 2252 33212
rect 1956 33158 2002 33210
rect 2002 33158 2012 33210
rect 2036 33158 2066 33210
rect 2066 33158 2078 33210
rect 2078 33158 2092 33210
rect 2116 33158 2130 33210
rect 2130 33158 2142 33210
rect 2142 33158 2172 33210
rect 2196 33158 2206 33210
rect 2206 33158 2252 33210
rect 1956 33156 2012 33158
rect 2036 33156 2092 33158
rect 2116 33156 2172 33158
rect 2196 33156 2252 33158
rect 6956 33210 7012 33212
rect 7036 33210 7092 33212
rect 7116 33210 7172 33212
rect 7196 33210 7252 33212
rect 6956 33158 7002 33210
rect 7002 33158 7012 33210
rect 7036 33158 7066 33210
rect 7066 33158 7078 33210
rect 7078 33158 7092 33210
rect 7116 33158 7130 33210
rect 7130 33158 7142 33210
rect 7142 33158 7172 33210
rect 7196 33158 7206 33210
rect 7206 33158 7252 33210
rect 6956 33156 7012 33158
rect 7036 33156 7092 33158
rect 7116 33156 7172 33158
rect 7196 33156 7252 33158
rect 11956 33210 12012 33212
rect 12036 33210 12092 33212
rect 12116 33210 12172 33212
rect 12196 33210 12252 33212
rect 11956 33158 12002 33210
rect 12002 33158 12012 33210
rect 12036 33158 12066 33210
rect 12066 33158 12078 33210
rect 12078 33158 12092 33210
rect 12116 33158 12130 33210
rect 12130 33158 12142 33210
rect 12142 33158 12172 33210
rect 12196 33158 12206 33210
rect 12206 33158 12252 33210
rect 11956 33156 12012 33158
rect 12036 33156 12092 33158
rect 12116 33156 12172 33158
rect 12196 33156 12252 33158
rect 16956 33210 17012 33212
rect 17036 33210 17092 33212
rect 17116 33210 17172 33212
rect 17196 33210 17252 33212
rect 16956 33158 17002 33210
rect 17002 33158 17012 33210
rect 17036 33158 17066 33210
rect 17066 33158 17078 33210
rect 17078 33158 17092 33210
rect 17116 33158 17130 33210
rect 17130 33158 17142 33210
rect 17142 33158 17172 33210
rect 17196 33158 17206 33210
rect 17206 33158 17252 33210
rect 16956 33156 17012 33158
rect 17036 33156 17092 33158
rect 17116 33156 17172 33158
rect 17196 33156 17252 33158
rect 21956 33210 22012 33212
rect 22036 33210 22092 33212
rect 22116 33210 22172 33212
rect 22196 33210 22252 33212
rect 21956 33158 22002 33210
rect 22002 33158 22012 33210
rect 22036 33158 22066 33210
rect 22066 33158 22078 33210
rect 22078 33158 22092 33210
rect 22116 33158 22130 33210
rect 22130 33158 22142 33210
rect 22142 33158 22172 33210
rect 22196 33158 22206 33210
rect 22206 33158 22252 33210
rect 21956 33156 22012 33158
rect 22036 33156 22092 33158
rect 22116 33156 22172 33158
rect 22196 33156 22252 33158
rect 26956 33210 27012 33212
rect 27036 33210 27092 33212
rect 27116 33210 27172 33212
rect 27196 33210 27252 33212
rect 26956 33158 27002 33210
rect 27002 33158 27012 33210
rect 27036 33158 27066 33210
rect 27066 33158 27078 33210
rect 27078 33158 27092 33210
rect 27116 33158 27130 33210
rect 27130 33158 27142 33210
rect 27142 33158 27172 33210
rect 27196 33158 27206 33210
rect 27206 33158 27252 33210
rect 26956 33156 27012 33158
rect 27036 33156 27092 33158
rect 27116 33156 27172 33158
rect 27196 33156 27252 33158
rect 31956 33210 32012 33212
rect 32036 33210 32092 33212
rect 32116 33210 32172 33212
rect 32196 33210 32252 33212
rect 31956 33158 32002 33210
rect 32002 33158 32012 33210
rect 32036 33158 32066 33210
rect 32066 33158 32078 33210
rect 32078 33158 32092 33210
rect 32116 33158 32130 33210
rect 32130 33158 32142 33210
rect 32142 33158 32172 33210
rect 32196 33158 32206 33210
rect 32206 33158 32252 33210
rect 31956 33156 32012 33158
rect 32036 33156 32092 33158
rect 32116 33156 32172 33158
rect 32196 33156 32252 33158
rect 36956 33210 37012 33212
rect 37036 33210 37092 33212
rect 37116 33210 37172 33212
rect 37196 33210 37252 33212
rect 36956 33158 37002 33210
rect 37002 33158 37012 33210
rect 37036 33158 37066 33210
rect 37066 33158 37078 33210
rect 37078 33158 37092 33210
rect 37116 33158 37130 33210
rect 37130 33158 37142 33210
rect 37142 33158 37172 33210
rect 37196 33158 37206 33210
rect 37206 33158 37252 33210
rect 36956 33156 37012 33158
rect 37036 33156 37092 33158
rect 37116 33156 37172 33158
rect 37196 33156 37252 33158
rect 2616 32666 2672 32668
rect 2696 32666 2752 32668
rect 2776 32666 2832 32668
rect 2856 32666 2912 32668
rect 2616 32614 2662 32666
rect 2662 32614 2672 32666
rect 2696 32614 2726 32666
rect 2726 32614 2738 32666
rect 2738 32614 2752 32666
rect 2776 32614 2790 32666
rect 2790 32614 2802 32666
rect 2802 32614 2832 32666
rect 2856 32614 2866 32666
rect 2866 32614 2912 32666
rect 2616 32612 2672 32614
rect 2696 32612 2752 32614
rect 2776 32612 2832 32614
rect 2856 32612 2912 32614
rect 7616 32666 7672 32668
rect 7696 32666 7752 32668
rect 7776 32666 7832 32668
rect 7856 32666 7912 32668
rect 7616 32614 7662 32666
rect 7662 32614 7672 32666
rect 7696 32614 7726 32666
rect 7726 32614 7738 32666
rect 7738 32614 7752 32666
rect 7776 32614 7790 32666
rect 7790 32614 7802 32666
rect 7802 32614 7832 32666
rect 7856 32614 7866 32666
rect 7866 32614 7912 32666
rect 7616 32612 7672 32614
rect 7696 32612 7752 32614
rect 7776 32612 7832 32614
rect 7856 32612 7912 32614
rect 12616 32666 12672 32668
rect 12696 32666 12752 32668
rect 12776 32666 12832 32668
rect 12856 32666 12912 32668
rect 12616 32614 12662 32666
rect 12662 32614 12672 32666
rect 12696 32614 12726 32666
rect 12726 32614 12738 32666
rect 12738 32614 12752 32666
rect 12776 32614 12790 32666
rect 12790 32614 12802 32666
rect 12802 32614 12832 32666
rect 12856 32614 12866 32666
rect 12866 32614 12912 32666
rect 12616 32612 12672 32614
rect 12696 32612 12752 32614
rect 12776 32612 12832 32614
rect 12856 32612 12912 32614
rect 17616 32666 17672 32668
rect 17696 32666 17752 32668
rect 17776 32666 17832 32668
rect 17856 32666 17912 32668
rect 17616 32614 17662 32666
rect 17662 32614 17672 32666
rect 17696 32614 17726 32666
rect 17726 32614 17738 32666
rect 17738 32614 17752 32666
rect 17776 32614 17790 32666
rect 17790 32614 17802 32666
rect 17802 32614 17832 32666
rect 17856 32614 17866 32666
rect 17866 32614 17912 32666
rect 17616 32612 17672 32614
rect 17696 32612 17752 32614
rect 17776 32612 17832 32614
rect 17856 32612 17912 32614
rect 22616 32666 22672 32668
rect 22696 32666 22752 32668
rect 22776 32666 22832 32668
rect 22856 32666 22912 32668
rect 22616 32614 22662 32666
rect 22662 32614 22672 32666
rect 22696 32614 22726 32666
rect 22726 32614 22738 32666
rect 22738 32614 22752 32666
rect 22776 32614 22790 32666
rect 22790 32614 22802 32666
rect 22802 32614 22832 32666
rect 22856 32614 22866 32666
rect 22866 32614 22912 32666
rect 22616 32612 22672 32614
rect 22696 32612 22752 32614
rect 22776 32612 22832 32614
rect 22856 32612 22912 32614
rect 27616 32666 27672 32668
rect 27696 32666 27752 32668
rect 27776 32666 27832 32668
rect 27856 32666 27912 32668
rect 27616 32614 27662 32666
rect 27662 32614 27672 32666
rect 27696 32614 27726 32666
rect 27726 32614 27738 32666
rect 27738 32614 27752 32666
rect 27776 32614 27790 32666
rect 27790 32614 27802 32666
rect 27802 32614 27832 32666
rect 27856 32614 27866 32666
rect 27866 32614 27912 32666
rect 27616 32612 27672 32614
rect 27696 32612 27752 32614
rect 27776 32612 27832 32614
rect 27856 32612 27912 32614
rect 32616 32666 32672 32668
rect 32696 32666 32752 32668
rect 32776 32666 32832 32668
rect 32856 32666 32912 32668
rect 32616 32614 32662 32666
rect 32662 32614 32672 32666
rect 32696 32614 32726 32666
rect 32726 32614 32738 32666
rect 32738 32614 32752 32666
rect 32776 32614 32790 32666
rect 32790 32614 32802 32666
rect 32802 32614 32832 32666
rect 32856 32614 32866 32666
rect 32866 32614 32912 32666
rect 32616 32612 32672 32614
rect 32696 32612 32752 32614
rect 32776 32612 32832 32614
rect 32856 32612 32912 32614
rect 37616 32666 37672 32668
rect 37696 32666 37752 32668
rect 37776 32666 37832 32668
rect 37856 32666 37912 32668
rect 37616 32614 37662 32666
rect 37662 32614 37672 32666
rect 37696 32614 37726 32666
rect 37726 32614 37738 32666
rect 37738 32614 37752 32666
rect 37776 32614 37790 32666
rect 37790 32614 37802 32666
rect 37802 32614 37832 32666
rect 37856 32614 37866 32666
rect 37866 32614 37912 32666
rect 37616 32612 37672 32614
rect 37696 32612 37752 32614
rect 37776 32612 37832 32614
rect 37856 32612 37912 32614
rect 1956 32122 2012 32124
rect 2036 32122 2092 32124
rect 2116 32122 2172 32124
rect 2196 32122 2252 32124
rect 1956 32070 2002 32122
rect 2002 32070 2012 32122
rect 2036 32070 2066 32122
rect 2066 32070 2078 32122
rect 2078 32070 2092 32122
rect 2116 32070 2130 32122
rect 2130 32070 2142 32122
rect 2142 32070 2172 32122
rect 2196 32070 2206 32122
rect 2206 32070 2252 32122
rect 1956 32068 2012 32070
rect 2036 32068 2092 32070
rect 2116 32068 2172 32070
rect 2196 32068 2252 32070
rect 6956 32122 7012 32124
rect 7036 32122 7092 32124
rect 7116 32122 7172 32124
rect 7196 32122 7252 32124
rect 6956 32070 7002 32122
rect 7002 32070 7012 32122
rect 7036 32070 7066 32122
rect 7066 32070 7078 32122
rect 7078 32070 7092 32122
rect 7116 32070 7130 32122
rect 7130 32070 7142 32122
rect 7142 32070 7172 32122
rect 7196 32070 7206 32122
rect 7206 32070 7252 32122
rect 6956 32068 7012 32070
rect 7036 32068 7092 32070
rect 7116 32068 7172 32070
rect 7196 32068 7252 32070
rect 11956 32122 12012 32124
rect 12036 32122 12092 32124
rect 12116 32122 12172 32124
rect 12196 32122 12252 32124
rect 11956 32070 12002 32122
rect 12002 32070 12012 32122
rect 12036 32070 12066 32122
rect 12066 32070 12078 32122
rect 12078 32070 12092 32122
rect 12116 32070 12130 32122
rect 12130 32070 12142 32122
rect 12142 32070 12172 32122
rect 12196 32070 12206 32122
rect 12206 32070 12252 32122
rect 11956 32068 12012 32070
rect 12036 32068 12092 32070
rect 12116 32068 12172 32070
rect 12196 32068 12252 32070
rect 16956 32122 17012 32124
rect 17036 32122 17092 32124
rect 17116 32122 17172 32124
rect 17196 32122 17252 32124
rect 16956 32070 17002 32122
rect 17002 32070 17012 32122
rect 17036 32070 17066 32122
rect 17066 32070 17078 32122
rect 17078 32070 17092 32122
rect 17116 32070 17130 32122
rect 17130 32070 17142 32122
rect 17142 32070 17172 32122
rect 17196 32070 17206 32122
rect 17206 32070 17252 32122
rect 16956 32068 17012 32070
rect 17036 32068 17092 32070
rect 17116 32068 17172 32070
rect 17196 32068 17252 32070
rect 21956 32122 22012 32124
rect 22036 32122 22092 32124
rect 22116 32122 22172 32124
rect 22196 32122 22252 32124
rect 21956 32070 22002 32122
rect 22002 32070 22012 32122
rect 22036 32070 22066 32122
rect 22066 32070 22078 32122
rect 22078 32070 22092 32122
rect 22116 32070 22130 32122
rect 22130 32070 22142 32122
rect 22142 32070 22172 32122
rect 22196 32070 22206 32122
rect 22206 32070 22252 32122
rect 21956 32068 22012 32070
rect 22036 32068 22092 32070
rect 22116 32068 22172 32070
rect 22196 32068 22252 32070
rect 26956 32122 27012 32124
rect 27036 32122 27092 32124
rect 27116 32122 27172 32124
rect 27196 32122 27252 32124
rect 26956 32070 27002 32122
rect 27002 32070 27012 32122
rect 27036 32070 27066 32122
rect 27066 32070 27078 32122
rect 27078 32070 27092 32122
rect 27116 32070 27130 32122
rect 27130 32070 27142 32122
rect 27142 32070 27172 32122
rect 27196 32070 27206 32122
rect 27206 32070 27252 32122
rect 26956 32068 27012 32070
rect 27036 32068 27092 32070
rect 27116 32068 27172 32070
rect 27196 32068 27252 32070
rect 31956 32122 32012 32124
rect 32036 32122 32092 32124
rect 32116 32122 32172 32124
rect 32196 32122 32252 32124
rect 31956 32070 32002 32122
rect 32002 32070 32012 32122
rect 32036 32070 32066 32122
rect 32066 32070 32078 32122
rect 32078 32070 32092 32122
rect 32116 32070 32130 32122
rect 32130 32070 32142 32122
rect 32142 32070 32172 32122
rect 32196 32070 32206 32122
rect 32206 32070 32252 32122
rect 31956 32068 32012 32070
rect 32036 32068 32092 32070
rect 32116 32068 32172 32070
rect 32196 32068 32252 32070
rect 36956 32122 37012 32124
rect 37036 32122 37092 32124
rect 37116 32122 37172 32124
rect 37196 32122 37252 32124
rect 36956 32070 37002 32122
rect 37002 32070 37012 32122
rect 37036 32070 37066 32122
rect 37066 32070 37078 32122
rect 37078 32070 37092 32122
rect 37116 32070 37130 32122
rect 37130 32070 37142 32122
rect 37142 32070 37172 32122
rect 37196 32070 37206 32122
rect 37206 32070 37252 32122
rect 36956 32068 37012 32070
rect 37036 32068 37092 32070
rect 37116 32068 37172 32070
rect 37196 32068 37252 32070
rect 2616 31578 2672 31580
rect 2696 31578 2752 31580
rect 2776 31578 2832 31580
rect 2856 31578 2912 31580
rect 2616 31526 2662 31578
rect 2662 31526 2672 31578
rect 2696 31526 2726 31578
rect 2726 31526 2738 31578
rect 2738 31526 2752 31578
rect 2776 31526 2790 31578
rect 2790 31526 2802 31578
rect 2802 31526 2832 31578
rect 2856 31526 2866 31578
rect 2866 31526 2912 31578
rect 2616 31524 2672 31526
rect 2696 31524 2752 31526
rect 2776 31524 2832 31526
rect 2856 31524 2912 31526
rect 7616 31578 7672 31580
rect 7696 31578 7752 31580
rect 7776 31578 7832 31580
rect 7856 31578 7912 31580
rect 7616 31526 7662 31578
rect 7662 31526 7672 31578
rect 7696 31526 7726 31578
rect 7726 31526 7738 31578
rect 7738 31526 7752 31578
rect 7776 31526 7790 31578
rect 7790 31526 7802 31578
rect 7802 31526 7832 31578
rect 7856 31526 7866 31578
rect 7866 31526 7912 31578
rect 7616 31524 7672 31526
rect 7696 31524 7752 31526
rect 7776 31524 7832 31526
rect 7856 31524 7912 31526
rect 12616 31578 12672 31580
rect 12696 31578 12752 31580
rect 12776 31578 12832 31580
rect 12856 31578 12912 31580
rect 12616 31526 12662 31578
rect 12662 31526 12672 31578
rect 12696 31526 12726 31578
rect 12726 31526 12738 31578
rect 12738 31526 12752 31578
rect 12776 31526 12790 31578
rect 12790 31526 12802 31578
rect 12802 31526 12832 31578
rect 12856 31526 12866 31578
rect 12866 31526 12912 31578
rect 12616 31524 12672 31526
rect 12696 31524 12752 31526
rect 12776 31524 12832 31526
rect 12856 31524 12912 31526
rect 17616 31578 17672 31580
rect 17696 31578 17752 31580
rect 17776 31578 17832 31580
rect 17856 31578 17912 31580
rect 17616 31526 17662 31578
rect 17662 31526 17672 31578
rect 17696 31526 17726 31578
rect 17726 31526 17738 31578
rect 17738 31526 17752 31578
rect 17776 31526 17790 31578
rect 17790 31526 17802 31578
rect 17802 31526 17832 31578
rect 17856 31526 17866 31578
rect 17866 31526 17912 31578
rect 17616 31524 17672 31526
rect 17696 31524 17752 31526
rect 17776 31524 17832 31526
rect 17856 31524 17912 31526
rect 22616 31578 22672 31580
rect 22696 31578 22752 31580
rect 22776 31578 22832 31580
rect 22856 31578 22912 31580
rect 22616 31526 22662 31578
rect 22662 31526 22672 31578
rect 22696 31526 22726 31578
rect 22726 31526 22738 31578
rect 22738 31526 22752 31578
rect 22776 31526 22790 31578
rect 22790 31526 22802 31578
rect 22802 31526 22832 31578
rect 22856 31526 22866 31578
rect 22866 31526 22912 31578
rect 22616 31524 22672 31526
rect 22696 31524 22752 31526
rect 22776 31524 22832 31526
rect 22856 31524 22912 31526
rect 27616 31578 27672 31580
rect 27696 31578 27752 31580
rect 27776 31578 27832 31580
rect 27856 31578 27912 31580
rect 27616 31526 27662 31578
rect 27662 31526 27672 31578
rect 27696 31526 27726 31578
rect 27726 31526 27738 31578
rect 27738 31526 27752 31578
rect 27776 31526 27790 31578
rect 27790 31526 27802 31578
rect 27802 31526 27832 31578
rect 27856 31526 27866 31578
rect 27866 31526 27912 31578
rect 27616 31524 27672 31526
rect 27696 31524 27752 31526
rect 27776 31524 27832 31526
rect 27856 31524 27912 31526
rect 32616 31578 32672 31580
rect 32696 31578 32752 31580
rect 32776 31578 32832 31580
rect 32856 31578 32912 31580
rect 32616 31526 32662 31578
rect 32662 31526 32672 31578
rect 32696 31526 32726 31578
rect 32726 31526 32738 31578
rect 32738 31526 32752 31578
rect 32776 31526 32790 31578
rect 32790 31526 32802 31578
rect 32802 31526 32832 31578
rect 32856 31526 32866 31578
rect 32866 31526 32912 31578
rect 32616 31524 32672 31526
rect 32696 31524 32752 31526
rect 32776 31524 32832 31526
rect 32856 31524 32912 31526
rect 37616 31578 37672 31580
rect 37696 31578 37752 31580
rect 37776 31578 37832 31580
rect 37856 31578 37912 31580
rect 37616 31526 37662 31578
rect 37662 31526 37672 31578
rect 37696 31526 37726 31578
rect 37726 31526 37738 31578
rect 37738 31526 37752 31578
rect 37776 31526 37790 31578
rect 37790 31526 37802 31578
rect 37802 31526 37832 31578
rect 37856 31526 37866 31578
rect 37866 31526 37912 31578
rect 37616 31524 37672 31526
rect 37696 31524 37752 31526
rect 37776 31524 37832 31526
rect 37856 31524 37912 31526
rect 1956 31034 2012 31036
rect 2036 31034 2092 31036
rect 2116 31034 2172 31036
rect 2196 31034 2252 31036
rect 1956 30982 2002 31034
rect 2002 30982 2012 31034
rect 2036 30982 2066 31034
rect 2066 30982 2078 31034
rect 2078 30982 2092 31034
rect 2116 30982 2130 31034
rect 2130 30982 2142 31034
rect 2142 30982 2172 31034
rect 2196 30982 2206 31034
rect 2206 30982 2252 31034
rect 1956 30980 2012 30982
rect 2036 30980 2092 30982
rect 2116 30980 2172 30982
rect 2196 30980 2252 30982
rect 6956 31034 7012 31036
rect 7036 31034 7092 31036
rect 7116 31034 7172 31036
rect 7196 31034 7252 31036
rect 6956 30982 7002 31034
rect 7002 30982 7012 31034
rect 7036 30982 7066 31034
rect 7066 30982 7078 31034
rect 7078 30982 7092 31034
rect 7116 30982 7130 31034
rect 7130 30982 7142 31034
rect 7142 30982 7172 31034
rect 7196 30982 7206 31034
rect 7206 30982 7252 31034
rect 6956 30980 7012 30982
rect 7036 30980 7092 30982
rect 7116 30980 7172 30982
rect 7196 30980 7252 30982
rect 11956 31034 12012 31036
rect 12036 31034 12092 31036
rect 12116 31034 12172 31036
rect 12196 31034 12252 31036
rect 11956 30982 12002 31034
rect 12002 30982 12012 31034
rect 12036 30982 12066 31034
rect 12066 30982 12078 31034
rect 12078 30982 12092 31034
rect 12116 30982 12130 31034
rect 12130 30982 12142 31034
rect 12142 30982 12172 31034
rect 12196 30982 12206 31034
rect 12206 30982 12252 31034
rect 11956 30980 12012 30982
rect 12036 30980 12092 30982
rect 12116 30980 12172 30982
rect 12196 30980 12252 30982
rect 16956 31034 17012 31036
rect 17036 31034 17092 31036
rect 17116 31034 17172 31036
rect 17196 31034 17252 31036
rect 16956 30982 17002 31034
rect 17002 30982 17012 31034
rect 17036 30982 17066 31034
rect 17066 30982 17078 31034
rect 17078 30982 17092 31034
rect 17116 30982 17130 31034
rect 17130 30982 17142 31034
rect 17142 30982 17172 31034
rect 17196 30982 17206 31034
rect 17206 30982 17252 31034
rect 16956 30980 17012 30982
rect 17036 30980 17092 30982
rect 17116 30980 17172 30982
rect 17196 30980 17252 30982
rect 21956 31034 22012 31036
rect 22036 31034 22092 31036
rect 22116 31034 22172 31036
rect 22196 31034 22252 31036
rect 21956 30982 22002 31034
rect 22002 30982 22012 31034
rect 22036 30982 22066 31034
rect 22066 30982 22078 31034
rect 22078 30982 22092 31034
rect 22116 30982 22130 31034
rect 22130 30982 22142 31034
rect 22142 30982 22172 31034
rect 22196 30982 22206 31034
rect 22206 30982 22252 31034
rect 21956 30980 22012 30982
rect 22036 30980 22092 30982
rect 22116 30980 22172 30982
rect 22196 30980 22252 30982
rect 26956 31034 27012 31036
rect 27036 31034 27092 31036
rect 27116 31034 27172 31036
rect 27196 31034 27252 31036
rect 26956 30982 27002 31034
rect 27002 30982 27012 31034
rect 27036 30982 27066 31034
rect 27066 30982 27078 31034
rect 27078 30982 27092 31034
rect 27116 30982 27130 31034
rect 27130 30982 27142 31034
rect 27142 30982 27172 31034
rect 27196 30982 27206 31034
rect 27206 30982 27252 31034
rect 26956 30980 27012 30982
rect 27036 30980 27092 30982
rect 27116 30980 27172 30982
rect 27196 30980 27252 30982
rect 31956 31034 32012 31036
rect 32036 31034 32092 31036
rect 32116 31034 32172 31036
rect 32196 31034 32252 31036
rect 31956 30982 32002 31034
rect 32002 30982 32012 31034
rect 32036 30982 32066 31034
rect 32066 30982 32078 31034
rect 32078 30982 32092 31034
rect 32116 30982 32130 31034
rect 32130 30982 32142 31034
rect 32142 30982 32172 31034
rect 32196 30982 32206 31034
rect 32206 30982 32252 31034
rect 31956 30980 32012 30982
rect 32036 30980 32092 30982
rect 32116 30980 32172 30982
rect 32196 30980 32252 30982
rect 36956 31034 37012 31036
rect 37036 31034 37092 31036
rect 37116 31034 37172 31036
rect 37196 31034 37252 31036
rect 36956 30982 37002 31034
rect 37002 30982 37012 31034
rect 37036 30982 37066 31034
rect 37066 30982 37078 31034
rect 37078 30982 37092 31034
rect 37116 30982 37130 31034
rect 37130 30982 37142 31034
rect 37142 30982 37172 31034
rect 37196 30982 37206 31034
rect 37206 30982 37252 31034
rect 36956 30980 37012 30982
rect 37036 30980 37092 30982
rect 37116 30980 37172 30982
rect 37196 30980 37252 30982
rect 2616 30490 2672 30492
rect 2696 30490 2752 30492
rect 2776 30490 2832 30492
rect 2856 30490 2912 30492
rect 2616 30438 2662 30490
rect 2662 30438 2672 30490
rect 2696 30438 2726 30490
rect 2726 30438 2738 30490
rect 2738 30438 2752 30490
rect 2776 30438 2790 30490
rect 2790 30438 2802 30490
rect 2802 30438 2832 30490
rect 2856 30438 2866 30490
rect 2866 30438 2912 30490
rect 2616 30436 2672 30438
rect 2696 30436 2752 30438
rect 2776 30436 2832 30438
rect 2856 30436 2912 30438
rect 7616 30490 7672 30492
rect 7696 30490 7752 30492
rect 7776 30490 7832 30492
rect 7856 30490 7912 30492
rect 7616 30438 7662 30490
rect 7662 30438 7672 30490
rect 7696 30438 7726 30490
rect 7726 30438 7738 30490
rect 7738 30438 7752 30490
rect 7776 30438 7790 30490
rect 7790 30438 7802 30490
rect 7802 30438 7832 30490
rect 7856 30438 7866 30490
rect 7866 30438 7912 30490
rect 7616 30436 7672 30438
rect 7696 30436 7752 30438
rect 7776 30436 7832 30438
rect 7856 30436 7912 30438
rect 12616 30490 12672 30492
rect 12696 30490 12752 30492
rect 12776 30490 12832 30492
rect 12856 30490 12912 30492
rect 12616 30438 12662 30490
rect 12662 30438 12672 30490
rect 12696 30438 12726 30490
rect 12726 30438 12738 30490
rect 12738 30438 12752 30490
rect 12776 30438 12790 30490
rect 12790 30438 12802 30490
rect 12802 30438 12832 30490
rect 12856 30438 12866 30490
rect 12866 30438 12912 30490
rect 12616 30436 12672 30438
rect 12696 30436 12752 30438
rect 12776 30436 12832 30438
rect 12856 30436 12912 30438
rect 17616 30490 17672 30492
rect 17696 30490 17752 30492
rect 17776 30490 17832 30492
rect 17856 30490 17912 30492
rect 17616 30438 17662 30490
rect 17662 30438 17672 30490
rect 17696 30438 17726 30490
rect 17726 30438 17738 30490
rect 17738 30438 17752 30490
rect 17776 30438 17790 30490
rect 17790 30438 17802 30490
rect 17802 30438 17832 30490
rect 17856 30438 17866 30490
rect 17866 30438 17912 30490
rect 17616 30436 17672 30438
rect 17696 30436 17752 30438
rect 17776 30436 17832 30438
rect 17856 30436 17912 30438
rect 22616 30490 22672 30492
rect 22696 30490 22752 30492
rect 22776 30490 22832 30492
rect 22856 30490 22912 30492
rect 22616 30438 22662 30490
rect 22662 30438 22672 30490
rect 22696 30438 22726 30490
rect 22726 30438 22738 30490
rect 22738 30438 22752 30490
rect 22776 30438 22790 30490
rect 22790 30438 22802 30490
rect 22802 30438 22832 30490
rect 22856 30438 22866 30490
rect 22866 30438 22912 30490
rect 22616 30436 22672 30438
rect 22696 30436 22752 30438
rect 22776 30436 22832 30438
rect 22856 30436 22912 30438
rect 27616 30490 27672 30492
rect 27696 30490 27752 30492
rect 27776 30490 27832 30492
rect 27856 30490 27912 30492
rect 27616 30438 27662 30490
rect 27662 30438 27672 30490
rect 27696 30438 27726 30490
rect 27726 30438 27738 30490
rect 27738 30438 27752 30490
rect 27776 30438 27790 30490
rect 27790 30438 27802 30490
rect 27802 30438 27832 30490
rect 27856 30438 27866 30490
rect 27866 30438 27912 30490
rect 27616 30436 27672 30438
rect 27696 30436 27752 30438
rect 27776 30436 27832 30438
rect 27856 30436 27912 30438
rect 32616 30490 32672 30492
rect 32696 30490 32752 30492
rect 32776 30490 32832 30492
rect 32856 30490 32912 30492
rect 32616 30438 32662 30490
rect 32662 30438 32672 30490
rect 32696 30438 32726 30490
rect 32726 30438 32738 30490
rect 32738 30438 32752 30490
rect 32776 30438 32790 30490
rect 32790 30438 32802 30490
rect 32802 30438 32832 30490
rect 32856 30438 32866 30490
rect 32866 30438 32912 30490
rect 32616 30436 32672 30438
rect 32696 30436 32752 30438
rect 32776 30436 32832 30438
rect 32856 30436 32912 30438
rect 37616 30490 37672 30492
rect 37696 30490 37752 30492
rect 37776 30490 37832 30492
rect 37856 30490 37912 30492
rect 37616 30438 37662 30490
rect 37662 30438 37672 30490
rect 37696 30438 37726 30490
rect 37726 30438 37738 30490
rect 37738 30438 37752 30490
rect 37776 30438 37790 30490
rect 37790 30438 37802 30490
rect 37802 30438 37832 30490
rect 37856 30438 37866 30490
rect 37866 30438 37912 30490
rect 37616 30436 37672 30438
rect 37696 30436 37752 30438
rect 37776 30436 37832 30438
rect 37856 30436 37912 30438
rect 1956 29946 2012 29948
rect 2036 29946 2092 29948
rect 2116 29946 2172 29948
rect 2196 29946 2252 29948
rect 1956 29894 2002 29946
rect 2002 29894 2012 29946
rect 2036 29894 2066 29946
rect 2066 29894 2078 29946
rect 2078 29894 2092 29946
rect 2116 29894 2130 29946
rect 2130 29894 2142 29946
rect 2142 29894 2172 29946
rect 2196 29894 2206 29946
rect 2206 29894 2252 29946
rect 1956 29892 2012 29894
rect 2036 29892 2092 29894
rect 2116 29892 2172 29894
rect 2196 29892 2252 29894
rect 6956 29946 7012 29948
rect 7036 29946 7092 29948
rect 7116 29946 7172 29948
rect 7196 29946 7252 29948
rect 6956 29894 7002 29946
rect 7002 29894 7012 29946
rect 7036 29894 7066 29946
rect 7066 29894 7078 29946
rect 7078 29894 7092 29946
rect 7116 29894 7130 29946
rect 7130 29894 7142 29946
rect 7142 29894 7172 29946
rect 7196 29894 7206 29946
rect 7206 29894 7252 29946
rect 6956 29892 7012 29894
rect 7036 29892 7092 29894
rect 7116 29892 7172 29894
rect 7196 29892 7252 29894
rect 11956 29946 12012 29948
rect 12036 29946 12092 29948
rect 12116 29946 12172 29948
rect 12196 29946 12252 29948
rect 11956 29894 12002 29946
rect 12002 29894 12012 29946
rect 12036 29894 12066 29946
rect 12066 29894 12078 29946
rect 12078 29894 12092 29946
rect 12116 29894 12130 29946
rect 12130 29894 12142 29946
rect 12142 29894 12172 29946
rect 12196 29894 12206 29946
rect 12206 29894 12252 29946
rect 11956 29892 12012 29894
rect 12036 29892 12092 29894
rect 12116 29892 12172 29894
rect 12196 29892 12252 29894
rect 16956 29946 17012 29948
rect 17036 29946 17092 29948
rect 17116 29946 17172 29948
rect 17196 29946 17252 29948
rect 16956 29894 17002 29946
rect 17002 29894 17012 29946
rect 17036 29894 17066 29946
rect 17066 29894 17078 29946
rect 17078 29894 17092 29946
rect 17116 29894 17130 29946
rect 17130 29894 17142 29946
rect 17142 29894 17172 29946
rect 17196 29894 17206 29946
rect 17206 29894 17252 29946
rect 16956 29892 17012 29894
rect 17036 29892 17092 29894
rect 17116 29892 17172 29894
rect 17196 29892 17252 29894
rect 21956 29946 22012 29948
rect 22036 29946 22092 29948
rect 22116 29946 22172 29948
rect 22196 29946 22252 29948
rect 21956 29894 22002 29946
rect 22002 29894 22012 29946
rect 22036 29894 22066 29946
rect 22066 29894 22078 29946
rect 22078 29894 22092 29946
rect 22116 29894 22130 29946
rect 22130 29894 22142 29946
rect 22142 29894 22172 29946
rect 22196 29894 22206 29946
rect 22206 29894 22252 29946
rect 21956 29892 22012 29894
rect 22036 29892 22092 29894
rect 22116 29892 22172 29894
rect 22196 29892 22252 29894
rect 26956 29946 27012 29948
rect 27036 29946 27092 29948
rect 27116 29946 27172 29948
rect 27196 29946 27252 29948
rect 26956 29894 27002 29946
rect 27002 29894 27012 29946
rect 27036 29894 27066 29946
rect 27066 29894 27078 29946
rect 27078 29894 27092 29946
rect 27116 29894 27130 29946
rect 27130 29894 27142 29946
rect 27142 29894 27172 29946
rect 27196 29894 27206 29946
rect 27206 29894 27252 29946
rect 26956 29892 27012 29894
rect 27036 29892 27092 29894
rect 27116 29892 27172 29894
rect 27196 29892 27252 29894
rect 31956 29946 32012 29948
rect 32036 29946 32092 29948
rect 32116 29946 32172 29948
rect 32196 29946 32252 29948
rect 31956 29894 32002 29946
rect 32002 29894 32012 29946
rect 32036 29894 32066 29946
rect 32066 29894 32078 29946
rect 32078 29894 32092 29946
rect 32116 29894 32130 29946
rect 32130 29894 32142 29946
rect 32142 29894 32172 29946
rect 32196 29894 32206 29946
rect 32206 29894 32252 29946
rect 31956 29892 32012 29894
rect 32036 29892 32092 29894
rect 32116 29892 32172 29894
rect 32196 29892 32252 29894
rect 36956 29946 37012 29948
rect 37036 29946 37092 29948
rect 37116 29946 37172 29948
rect 37196 29946 37252 29948
rect 36956 29894 37002 29946
rect 37002 29894 37012 29946
rect 37036 29894 37066 29946
rect 37066 29894 37078 29946
rect 37078 29894 37092 29946
rect 37116 29894 37130 29946
rect 37130 29894 37142 29946
rect 37142 29894 37172 29946
rect 37196 29894 37206 29946
rect 37206 29894 37252 29946
rect 36956 29892 37012 29894
rect 37036 29892 37092 29894
rect 37116 29892 37172 29894
rect 37196 29892 37252 29894
rect 2616 29402 2672 29404
rect 2696 29402 2752 29404
rect 2776 29402 2832 29404
rect 2856 29402 2912 29404
rect 2616 29350 2662 29402
rect 2662 29350 2672 29402
rect 2696 29350 2726 29402
rect 2726 29350 2738 29402
rect 2738 29350 2752 29402
rect 2776 29350 2790 29402
rect 2790 29350 2802 29402
rect 2802 29350 2832 29402
rect 2856 29350 2866 29402
rect 2866 29350 2912 29402
rect 2616 29348 2672 29350
rect 2696 29348 2752 29350
rect 2776 29348 2832 29350
rect 2856 29348 2912 29350
rect 7616 29402 7672 29404
rect 7696 29402 7752 29404
rect 7776 29402 7832 29404
rect 7856 29402 7912 29404
rect 7616 29350 7662 29402
rect 7662 29350 7672 29402
rect 7696 29350 7726 29402
rect 7726 29350 7738 29402
rect 7738 29350 7752 29402
rect 7776 29350 7790 29402
rect 7790 29350 7802 29402
rect 7802 29350 7832 29402
rect 7856 29350 7866 29402
rect 7866 29350 7912 29402
rect 7616 29348 7672 29350
rect 7696 29348 7752 29350
rect 7776 29348 7832 29350
rect 7856 29348 7912 29350
rect 12616 29402 12672 29404
rect 12696 29402 12752 29404
rect 12776 29402 12832 29404
rect 12856 29402 12912 29404
rect 12616 29350 12662 29402
rect 12662 29350 12672 29402
rect 12696 29350 12726 29402
rect 12726 29350 12738 29402
rect 12738 29350 12752 29402
rect 12776 29350 12790 29402
rect 12790 29350 12802 29402
rect 12802 29350 12832 29402
rect 12856 29350 12866 29402
rect 12866 29350 12912 29402
rect 12616 29348 12672 29350
rect 12696 29348 12752 29350
rect 12776 29348 12832 29350
rect 12856 29348 12912 29350
rect 17616 29402 17672 29404
rect 17696 29402 17752 29404
rect 17776 29402 17832 29404
rect 17856 29402 17912 29404
rect 17616 29350 17662 29402
rect 17662 29350 17672 29402
rect 17696 29350 17726 29402
rect 17726 29350 17738 29402
rect 17738 29350 17752 29402
rect 17776 29350 17790 29402
rect 17790 29350 17802 29402
rect 17802 29350 17832 29402
rect 17856 29350 17866 29402
rect 17866 29350 17912 29402
rect 17616 29348 17672 29350
rect 17696 29348 17752 29350
rect 17776 29348 17832 29350
rect 17856 29348 17912 29350
rect 22616 29402 22672 29404
rect 22696 29402 22752 29404
rect 22776 29402 22832 29404
rect 22856 29402 22912 29404
rect 22616 29350 22662 29402
rect 22662 29350 22672 29402
rect 22696 29350 22726 29402
rect 22726 29350 22738 29402
rect 22738 29350 22752 29402
rect 22776 29350 22790 29402
rect 22790 29350 22802 29402
rect 22802 29350 22832 29402
rect 22856 29350 22866 29402
rect 22866 29350 22912 29402
rect 22616 29348 22672 29350
rect 22696 29348 22752 29350
rect 22776 29348 22832 29350
rect 22856 29348 22912 29350
rect 27616 29402 27672 29404
rect 27696 29402 27752 29404
rect 27776 29402 27832 29404
rect 27856 29402 27912 29404
rect 27616 29350 27662 29402
rect 27662 29350 27672 29402
rect 27696 29350 27726 29402
rect 27726 29350 27738 29402
rect 27738 29350 27752 29402
rect 27776 29350 27790 29402
rect 27790 29350 27802 29402
rect 27802 29350 27832 29402
rect 27856 29350 27866 29402
rect 27866 29350 27912 29402
rect 27616 29348 27672 29350
rect 27696 29348 27752 29350
rect 27776 29348 27832 29350
rect 27856 29348 27912 29350
rect 32616 29402 32672 29404
rect 32696 29402 32752 29404
rect 32776 29402 32832 29404
rect 32856 29402 32912 29404
rect 32616 29350 32662 29402
rect 32662 29350 32672 29402
rect 32696 29350 32726 29402
rect 32726 29350 32738 29402
rect 32738 29350 32752 29402
rect 32776 29350 32790 29402
rect 32790 29350 32802 29402
rect 32802 29350 32832 29402
rect 32856 29350 32866 29402
rect 32866 29350 32912 29402
rect 32616 29348 32672 29350
rect 32696 29348 32752 29350
rect 32776 29348 32832 29350
rect 32856 29348 32912 29350
rect 37616 29402 37672 29404
rect 37696 29402 37752 29404
rect 37776 29402 37832 29404
rect 37856 29402 37912 29404
rect 37616 29350 37662 29402
rect 37662 29350 37672 29402
rect 37696 29350 37726 29402
rect 37726 29350 37738 29402
rect 37738 29350 37752 29402
rect 37776 29350 37790 29402
rect 37790 29350 37802 29402
rect 37802 29350 37832 29402
rect 37856 29350 37866 29402
rect 37866 29350 37912 29402
rect 37616 29348 37672 29350
rect 37696 29348 37752 29350
rect 37776 29348 37832 29350
rect 37856 29348 37912 29350
rect 1956 28858 2012 28860
rect 2036 28858 2092 28860
rect 2116 28858 2172 28860
rect 2196 28858 2252 28860
rect 1956 28806 2002 28858
rect 2002 28806 2012 28858
rect 2036 28806 2066 28858
rect 2066 28806 2078 28858
rect 2078 28806 2092 28858
rect 2116 28806 2130 28858
rect 2130 28806 2142 28858
rect 2142 28806 2172 28858
rect 2196 28806 2206 28858
rect 2206 28806 2252 28858
rect 1956 28804 2012 28806
rect 2036 28804 2092 28806
rect 2116 28804 2172 28806
rect 2196 28804 2252 28806
rect 6956 28858 7012 28860
rect 7036 28858 7092 28860
rect 7116 28858 7172 28860
rect 7196 28858 7252 28860
rect 6956 28806 7002 28858
rect 7002 28806 7012 28858
rect 7036 28806 7066 28858
rect 7066 28806 7078 28858
rect 7078 28806 7092 28858
rect 7116 28806 7130 28858
rect 7130 28806 7142 28858
rect 7142 28806 7172 28858
rect 7196 28806 7206 28858
rect 7206 28806 7252 28858
rect 6956 28804 7012 28806
rect 7036 28804 7092 28806
rect 7116 28804 7172 28806
rect 7196 28804 7252 28806
rect 11956 28858 12012 28860
rect 12036 28858 12092 28860
rect 12116 28858 12172 28860
rect 12196 28858 12252 28860
rect 11956 28806 12002 28858
rect 12002 28806 12012 28858
rect 12036 28806 12066 28858
rect 12066 28806 12078 28858
rect 12078 28806 12092 28858
rect 12116 28806 12130 28858
rect 12130 28806 12142 28858
rect 12142 28806 12172 28858
rect 12196 28806 12206 28858
rect 12206 28806 12252 28858
rect 11956 28804 12012 28806
rect 12036 28804 12092 28806
rect 12116 28804 12172 28806
rect 12196 28804 12252 28806
rect 16956 28858 17012 28860
rect 17036 28858 17092 28860
rect 17116 28858 17172 28860
rect 17196 28858 17252 28860
rect 16956 28806 17002 28858
rect 17002 28806 17012 28858
rect 17036 28806 17066 28858
rect 17066 28806 17078 28858
rect 17078 28806 17092 28858
rect 17116 28806 17130 28858
rect 17130 28806 17142 28858
rect 17142 28806 17172 28858
rect 17196 28806 17206 28858
rect 17206 28806 17252 28858
rect 16956 28804 17012 28806
rect 17036 28804 17092 28806
rect 17116 28804 17172 28806
rect 17196 28804 17252 28806
rect 21956 28858 22012 28860
rect 22036 28858 22092 28860
rect 22116 28858 22172 28860
rect 22196 28858 22252 28860
rect 21956 28806 22002 28858
rect 22002 28806 22012 28858
rect 22036 28806 22066 28858
rect 22066 28806 22078 28858
rect 22078 28806 22092 28858
rect 22116 28806 22130 28858
rect 22130 28806 22142 28858
rect 22142 28806 22172 28858
rect 22196 28806 22206 28858
rect 22206 28806 22252 28858
rect 21956 28804 22012 28806
rect 22036 28804 22092 28806
rect 22116 28804 22172 28806
rect 22196 28804 22252 28806
rect 26956 28858 27012 28860
rect 27036 28858 27092 28860
rect 27116 28858 27172 28860
rect 27196 28858 27252 28860
rect 26956 28806 27002 28858
rect 27002 28806 27012 28858
rect 27036 28806 27066 28858
rect 27066 28806 27078 28858
rect 27078 28806 27092 28858
rect 27116 28806 27130 28858
rect 27130 28806 27142 28858
rect 27142 28806 27172 28858
rect 27196 28806 27206 28858
rect 27206 28806 27252 28858
rect 26956 28804 27012 28806
rect 27036 28804 27092 28806
rect 27116 28804 27172 28806
rect 27196 28804 27252 28806
rect 31956 28858 32012 28860
rect 32036 28858 32092 28860
rect 32116 28858 32172 28860
rect 32196 28858 32252 28860
rect 31956 28806 32002 28858
rect 32002 28806 32012 28858
rect 32036 28806 32066 28858
rect 32066 28806 32078 28858
rect 32078 28806 32092 28858
rect 32116 28806 32130 28858
rect 32130 28806 32142 28858
rect 32142 28806 32172 28858
rect 32196 28806 32206 28858
rect 32206 28806 32252 28858
rect 31956 28804 32012 28806
rect 32036 28804 32092 28806
rect 32116 28804 32172 28806
rect 32196 28804 32252 28806
rect 36956 28858 37012 28860
rect 37036 28858 37092 28860
rect 37116 28858 37172 28860
rect 37196 28858 37252 28860
rect 36956 28806 37002 28858
rect 37002 28806 37012 28858
rect 37036 28806 37066 28858
rect 37066 28806 37078 28858
rect 37078 28806 37092 28858
rect 37116 28806 37130 28858
rect 37130 28806 37142 28858
rect 37142 28806 37172 28858
rect 37196 28806 37206 28858
rect 37206 28806 37252 28858
rect 36956 28804 37012 28806
rect 37036 28804 37092 28806
rect 37116 28804 37172 28806
rect 37196 28804 37252 28806
rect 2616 28314 2672 28316
rect 2696 28314 2752 28316
rect 2776 28314 2832 28316
rect 2856 28314 2912 28316
rect 2616 28262 2662 28314
rect 2662 28262 2672 28314
rect 2696 28262 2726 28314
rect 2726 28262 2738 28314
rect 2738 28262 2752 28314
rect 2776 28262 2790 28314
rect 2790 28262 2802 28314
rect 2802 28262 2832 28314
rect 2856 28262 2866 28314
rect 2866 28262 2912 28314
rect 2616 28260 2672 28262
rect 2696 28260 2752 28262
rect 2776 28260 2832 28262
rect 2856 28260 2912 28262
rect 7616 28314 7672 28316
rect 7696 28314 7752 28316
rect 7776 28314 7832 28316
rect 7856 28314 7912 28316
rect 7616 28262 7662 28314
rect 7662 28262 7672 28314
rect 7696 28262 7726 28314
rect 7726 28262 7738 28314
rect 7738 28262 7752 28314
rect 7776 28262 7790 28314
rect 7790 28262 7802 28314
rect 7802 28262 7832 28314
rect 7856 28262 7866 28314
rect 7866 28262 7912 28314
rect 7616 28260 7672 28262
rect 7696 28260 7752 28262
rect 7776 28260 7832 28262
rect 7856 28260 7912 28262
rect 12616 28314 12672 28316
rect 12696 28314 12752 28316
rect 12776 28314 12832 28316
rect 12856 28314 12912 28316
rect 12616 28262 12662 28314
rect 12662 28262 12672 28314
rect 12696 28262 12726 28314
rect 12726 28262 12738 28314
rect 12738 28262 12752 28314
rect 12776 28262 12790 28314
rect 12790 28262 12802 28314
rect 12802 28262 12832 28314
rect 12856 28262 12866 28314
rect 12866 28262 12912 28314
rect 12616 28260 12672 28262
rect 12696 28260 12752 28262
rect 12776 28260 12832 28262
rect 12856 28260 12912 28262
rect 17616 28314 17672 28316
rect 17696 28314 17752 28316
rect 17776 28314 17832 28316
rect 17856 28314 17912 28316
rect 17616 28262 17662 28314
rect 17662 28262 17672 28314
rect 17696 28262 17726 28314
rect 17726 28262 17738 28314
rect 17738 28262 17752 28314
rect 17776 28262 17790 28314
rect 17790 28262 17802 28314
rect 17802 28262 17832 28314
rect 17856 28262 17866 28314
rect 17866 28262 17912 28314
rect 17616 28260 17672 28262
rect 17696 28260 17752 28262
rect 17776 28260 17832 28262
rect 17856 28260 17912 28262
rect 22616 28314 22672 28316
rect 22696 28314 22752 28316
rect 22776 28314 22832 28316
rect 22856 28314 22912 28316
rect 22616 28262 22662 28314
rect 22662 28262 22672 28314
rect 22696 28262 22726 28314
rect 22726 28262 22738 28314
rect 22738 28262 22752 28314
rect 22776 28262 22790 28314
rect 22790 28262 22802 28314
rect 22802 28262 22832 28314
rect 22856 28262 22866 28314
rect 22866 28262 22912 28314
rect 22616 28260 22672 28262
rect 22696 28260 22752 28262
rect 22776 28260 22832 28262
rect 22856 28260 22912 28262
rect 27616 28314 27672 28316
rect 27696 28314 27752 28316
rect 27776 28314 27832 28316
rect 27856 28314 27912 28316
rect 27616 28262 27662 28314
rect 27662 28262 27672 28314
rect 27696 28262 27726 28314
rect 27726 28262 27738 28314
rect 27738 28262 27752 28314
rect 27776 28262 27790 28314
rect 27790 28262 27802 28314
rect 27802 28262 27832 28314
rect 27856 28262 27866 28314
rect 27866 28262 27912 28314
rect 27616 28260 27672 28262
rect 27696 28260 27752 28262
rect 27776 28260 27832 28262
rect 27856 28260 27912 28262
rect 32616 28314 32672 28316
rect 32696 28314 32752 28316
rect 32776 28314 32832 28316
rect 32856 28314 32912 28316
rect 32616 28262 32662 28314
rect 32662 28262 32672 28314
rect 32696 28262 32726 28314
rect 32726 28262 32738 28314
rect 32738 28262 32752 28314
rect 32776 28262 32790 28314
rect 32790 28262 32802 28314
rect 32802 28262 32832 28314
rect 32856 28262 32866 28314
rect 32866 28262 32912 28314
rect 32616 28260 32672 28262
rect 32696 28260 32752 28262
rect 32776 28260 32832 28262
rect 32856 28260 32912 28262
rect 37616 28314 37672 28316
rect 37696 28314 37752 28316
rect 37776 28314 37832 28316
rect 37856 28314 37912 28316
rect 37616 28262 37662 28314
rect 37662 28262 37672 28314
rect 37696 28262 37726 28314
rect 37726 28262 37738 28314
rect 37738 28262 37752 28314
rect 37776 28262 37790 28314
rect 37790 28262 37802 28314
rect 37802 28262 37832 28314
rect 37856 28262 37866 28314
rect 37866 28262 37912 28314
rect 37616 28260 37672 28262
rect 37696 28260 37752 28262
rect 37776 28260 37832 28262
rect 37856 28260 37912 28262
rect 1956 27770 2012 27772
rect 2036 27770 2092 27772
rect 2116 27770 2172 27772
rect 2196 27770 2252 27772
rect 1956 27718 2002 27770
rect 2002 27718 2012 27770
rect 2036 27718 2066 27770
rect 2066 27718 2078 27770
rect 2078 27718 2092 27770
rect 2116 27718 2130 27770
rect 2130 27718 2142 27770
rect 2142 27718 2172 27770
rect 2196 27718 2206 27770
rect 2206 27718 2252 27770
rect 1956 27716 2012 27718
rect 2036 27716 2092 27718
rect 2116 27716 2172 27718
rect 2196 27716 2252 27718
rect 6956 27770 7012 27772
rect 7036 27770 7092 27772
rect 7116 27770 7172 27772
rect 7196 27770 7252 27772
rect 6956 27718 7002 27770
rect 7002 27718 7012 27770
rect 7036 27718 7066 27770
rect 7066 27718 7078 27770
rect 7078 27718 7092 27770
rect 7116 27718 7130 27770
rect 7130 27718 7142 27770
rect 7142 27718 7172 27770
rect 7196 27718 7206 27770
rect 7206 27718 7252 27770
rect 6956 27716 7012 27718
rect 7036 27716 7092 27718
rect 7116 27716 7172 27718
rect 7196 27716 7252 27718
rect 11956 27770 12012 27772
rect 12036 27770 12092 27772
rect 12116 27770 12172 27772
rect 12196 27770 12252 27772
rect 11956 27718 12002 27770
rect 12002 27718 12012 27770
rect 12036 27718 12066 27770
rect 12066 27718 12078 27770
rect 12078 27718 12092 27770
rect 12116 27718 12130 27770
rect 12130 27718 12142 27770
rect 12142 27718 12172 27770
rect 12196 27718 12206 27770
rect 12206 27718 12252 27770
rect 11956 27716 12012 27718
rect 12036 27716 12092 27718
rect 12116 27716 12172 27718
rect 12196 27716 12252 27718
rect 16956 27770 17012 27772
rect 17036 27770 17092 27772
rect 17116 27770 17172 27772
rect 17196 27770 17252 27772
rect 16956 27718 17002 27770
rect 17002 27718 17012 27770
rect 17036 27718 17066 27770
rect 17066 27718 17078 27770
rect 17078 27718 17092 27770
rect 17116 27718 17130 27770
rect 17130 27718 17142 27770
rect 17142 27718 17172 27770
rect 17196 27718 17206 27770
rect 17206 27718 17252 27770
rect 16956 27716 17012 27718
rect 17036 27716 17092 27718
rect 17116 27716 17172 27718
rect 17196 27716 17252 27718
rect 21956 27770 22012 27772
rect 22036 27770 22092 27772
rect 22116 27770 22172 27772
rect 22196 27770 22252 27772
rect 21956 27718 22002 27770
rect 22002 27718 22012 27770
rect 22036 27718 22066 27770
rect 22066 27718 22078 27770
rect 22078 27718 22092 27770
rect 22116 27718 22130 27770
rect 22130 27718 22142 27770
rect 22142 27718 22172 27770
rect 22196 27718 22206 27770
rect 22206 27718 22252 27770
rect 21956 27716 22012 27718
rect 22036 27716 22092 27718
rect 22116 27716 22172 27718
rect 22196 27716 22252 27718
rect 26956 27770 27012 27772
rect 27036 27770 27092 27772
rect 27116 27770 27172 27772
rect 27196 27770 27252 27772
rect 26956 27718 27002 27770
rect 27002 27718 27012 27770
rect 27036 27718 27066 27770
rect 27066 27718 27078 27770
rect 27078 27718 27092 27770
rect 27116 27718 27130 27770
rect 27130 27718 27142 27770
rect 27142 27718 27172 27770
rect 27196 27718 27206 27770
rect 27206 27718 27252 27770
rect 26956 27716 27012 27718
rect 27036 27716 27092 27718
rect 27116 27716 27172 27718
rect 27196 27716 27252 27718
rect 31956 27770 32012 27772
rect 32036 27770 32092 27772
rect 32116 27770 32172 27772
rect 32196 27770 32252 27772
rect 31956 27718 32002 27770
rect 32002 27718 32012 27770
rect 32036 27718 32066 27770
rect 32066 27718 32078 27770
rect 32078 27718 32092 27770
rect 32116 27718 32130 27770
rect 32130 27718 32142 27770
rect 32142 27718 32172 27770
rect 32196 27718 32206 27770
rect 32206 27718 32252 27770
rect 31956 27716 32012 27718
rect 32036 27716 32092 27718
rect 32116 27716 32172 27718
rect 32196 27716 32252 27718
rect 36956 27770 37012 27772
rect 37036 27770 37092 27772
rect 37116 27770 37172 27772
rect 37196 27770 37252 27772
rect 36956 27718 37002 27770
rect 37002 27718 37012 27770
rect 37036 27718 37066 27770
rect 37066 27718 37078 27770
rect 37078 27718 37092 27770
rect 37116 27718 37130 27770
rect 37130 27718 37142 27770
rect 37142 27718 37172 27770
rect 37196 27718 37206 27770
rect 37206 27718 37252 27770
rect 36956 27716 37012 27718
rect 37036 27716 37092 27718
rect 37116 27716 37172 27718
rect 37196 27716 37252 27718
rect 2616 27226 2672 27228
rect 2696 27226 2752 27228
rect 2776 27226 2832 27228
rect 2856 27226 2912 27228
rect 2616 27174 2662 27226
rect 2662 27174 2672 27226
rect 2696 27174 2726 27226
rect 2726 27174 2738 27226
rect 2738 27174 2752 27226
rect 2776 27174 2790 27226
rect 2790 27174 2802 27226
rect 2802 27174 2832 27226
rect 2856 27174 2866 27226
rect 2866 27174 2912 27226
rect 2616 27172 2672 27174
rect 2696 27172 2752 27174
rect 2776 27172 2832 27174
rect 2856 27172 2912 27174
rect 7616 27226 7672 27228
rect 7696 27226 7752 27228
rect 7776 27226 7832 27228
rect 7856 27226 7912 27228
rect 7616 27174 7662 27226
rect 7662 27174 7672 27226
rect 7696 27174 7726 27226
rect 7726 27174 7738 27226
rect 7738 27174 7752 27226
rect 7776 27174 7790 27226
rect 7790 27174 7802 27226
rect 7802 27174 7832 27226
rect 7856 27174 7866 27226
rect 7866 27174 7912 27226
rect 7616 27172 7672 27174
rect 7696 27172 7752 27174
rect 7776 27172 7832 27174
rect 7856 27172 7912 27174
rect 12616 27226 12672 27228
rect 12696 27226 12752 27228
rect 12776 27226 12832 27228
rect 12856 27226 12912 27228
rect 12616 27174 12662 27226
rect 12662 27174 12672 27226
rect 12696 27174 12726 27226
rect 12726 27174 12738 27226
rect 12738 27174 12752 27226
rect 12776 27174 12790 27226
rect 12790 27174 12802 27226
rect 12802 27174 12832 27226
rect 12856 27174 12866 27226
rect 12866 27174 12912 27226
rect 12616 27172 12672 27174
rect 12696 27172 12752 27174
rect 12776 27172 12832 27174
rect 12856 27172 12912 27174
rect 17616 27226 17672 27228
rect 17696 27226 17752 27228
rect 17776 27226 17832 27228
rect 17856 27226 17912 27228
rect 17616 27174 17662 27226
rect 17662 27174 17672 27226
rect 17696 27174 17726 27226
rect 17726 27174 17738 27226
rect 17738 27174 17752 27226
rect 17776 27174 17790 27226
rect 17790 27174 17802 27226
rect 17802 27174 17832 27226
rect 17856 27174 17866 27226
rect 17866 27174 17912 27226
rect 17616 27172 17672 27174
rect 17696 27172 17752 27174
rect 17776 27172 17832 27174
rect 17856 27172 17912 27174
rect 22616 27226 22672 27228
rect 22696 27226 22752 27228
rect 22776 27226 22832 27228
rect 22856 27226 22912 27228
rect 22616 27174 22662 27226
rect 22662 27174 22672 27226
rect 22696 27174 22726 27226
rect 22726 27174 22738 27226
rect 22738 27174 22752 27226
rect 22776 27174 22790 27226
rect 22790 27174 22802 27226
rect 22802 27174 22832 27226
rect 22856 27174 22866 27226
rect 22866 27174 22912 27226
rect 22616 27172 22672 27174
rect 22696 27172 22752 27174
rect 22776 27172 22832 27174
rect 22856 27172 22912 27174
rect 27616 27226 27672 27228
rect 27696 27226 27752 27228
rect 27776 27226 27832 27228
rect 27856 27226 27912 27228
rect 27616 27174 27662 27226
rect 27662 27174 27672 27226
rect 27696 27174 27726 27226
rect 27726 27174 27738 27226
rect 27738 27174 27752 27226
rect 27776 27174 27790 27226
rect 27790 27174 27802 27226
rect 27802 27174 27832 27226
rect 27856 27174 27866 27226
rect 27866 27174 27912 27226
rect 27616 27172 27672 27174
rect 27696 27172 27752 27174
rect 27776 27172 27832 27174
rect 27856 27172 27912 27174
rect 32616 27226 32672 27228
rect 32696 27226 32752 27228
rect 32776 27226 32832 27228
rect 32856 27226 32912 27228
rect 32616 27174 32662 27226
rect 32662 27174 32672 27226
rect 32696 27174 32726 27226
rect 32726 27174 32738 27226
rect 32738 27174 32752 27226
rect 32776 27174 32790 27226
rect 32790 27174 32802 27226
rect 32802 27174 32832 27226
rect 32856 27174 32866 27226
rect 32866 27174 32912 27226
rect 32616 27172 32672 27174
rect 32696 27172 32752 27174
rect 32776 27172 32832 27174
rect 32856 27172 32912 27174
rect 37616 27226 37672 27228
rect 37696 27226 37752 27228
rect 37776 27226 37832 27228
rect 37856 27226 37912 27228
rect 37616 27174 37662 27226
rect 37662 27174 37672 27226
rect 37696 27174 37726 27226
rect 37726 27174 37738 27226
rect 37738 27174 37752 27226
rect 37776 27174 37790 27226
rect 37790 27174 37802 27226
rect 37802 27174 37832 27226
rect 37856 27174 37866 27226
rect 37866 27174 37912 27226
rect 37616 27172 37672 27174
rect 37696 27172 37752 27174
rect 37776 27172 37832 27174
rect 37856 27172 37912 27174
rect 1956 26682 2012 26684
rect 2036 26682 2092 26684
rect 2116 26682 2172 26684
rect 2196 26682 2252 26684
rect 1956 26630 2002 26682
rect 2002 26630 2012 26682
rect 2036 26630 2066 26682
rect 2066 26630 2078 26682
rect 2078 26630 2092 26682
rect 2116 26630 2130 26682
rect 2130 26630 2142 26682
rect 2142 26630 2172 26682
rect 2196 26630 2206 26682
rect 2206 26630 2252 26682
rect 1956 26628 2012 26630
rect 2036 26628 2092 26630
rect 2116 26628 2172 26630
rect 2196 26628 2252 26630
rect 6956 26682 7012 26684
rect 7036 26682 7092 26684
rect 7116 26682 7172 26684
rect 7196 26682 7252 26684
rect 6956 26630 7002 26682
rect 7002 26630 7012 26682
rect 7036 26630 7066 26682
rect 7066 26630 7078 26682
rect 7078 26630 7092 26682
rect 7116 26630 7130 26682
rect 7130 26630 7142 26682
rect 7142 26630 7172 26682
rect 7196 26630 7206 26682
rect 7206 26630 7252 26682
rect 6956 26628 7012 26630
rect 7036 26628 7092 26630
rect 7116 26628 7172 26630
rect 7196 26628 7252 26630
rect 11956 26682 12012 26684
rect 12036 26682 12092 26684
rect 12116 26682 12172 26684
rect 12196 26682 12252 26684
rect 11956 26630 12002 26682
rect 12002 26630 12012 26682
rect 12036 26630 12066 26682
rect 12066 26630 12078 26682
rect 12078 26630 12092 26682
rect 12116 26630 12130 26682
rect 12130 26630 12142 26682
rect 12142 26630 12172 26682
rect 12196 26630 12206 26682
rect 12206 26630 12252 26682
rect 11956 26628 12012 26630
rect 12036 26628 12092 26630
rect 12116 26628 12172 26630
rect 12196 26628 12252 26630
rect 16956 26682 17012 26684
rect 17036 26682 17092 26684
rect 17116 26682 17172 26684
rect 17196 26682 17252 26684
rect 16956 26630 17002 26682
rect 17002 26630 17012 26682
rect 17036 26630 17066 26682
rect 17066 26630 17078 26682
rect 17078 26630 17092 26682
rect 17116 26630 17130 26682
rect 17130 26630 17142 26682
rect 17142 26630 17172 26682
rect 17196 26630 17206 26682
rect 17206 26630 17252 26682
rect 16956 26628 17012 26630
rect 17036 26628 17092 26630
rect 17116 26628 17172 26630
rect 17196 26628 17252 26630
rect 21956 26682 22012 26684
rect 22036 26682 22092 26684
rect 22116 26682 22172 26684
rect 22196 26682 22252 26684
rect 21956 26630 22002 26682
rect 22002 26630 22012 26682
rect 22036 26630 22066 26682
rect 22066 26630 22078 26682
rect 22078 26630 22092 26682
rect 22116 26630 22130 26682
rect 22130 26630 22142 26682
rect 22142 26630 22172 26682
rect 22196 26630 22206 26682
rect 22206 26630 22252 26682
rect 21956 26628 22012 26630
rect 22036 26628 22092 26630
rect 22116 26628 22172 26630
rect 22196 26628 22252 26630
rect 26956 26682 27012 26684
rect 27036 26682 27092 26684
rect 27116 26682 27172 26684
rect 27196 26682 27252 26684
rect 26956 26630 27002 26682
rect 27002 26630 27012 26682
rect 27036 26630 27066 26682
rect 27066 26630 27078 26682
rect 27078 26630 27092 26682
rect 27116 26630 27130 26682
rect 27130 26630 27142 26682
rect 27142 26630 27172 26682
rect 27196 26630 27206 26682
rect 27206 26630 27252 26682
rect 26956 26628 27012 26630
rect 27036 26628 27092 26630
rect 27116 26628 27172 26630
rect 27196 26628 27252 26630
rect 31956 26682 32012 26684
rect 32036 26682 32092 26684
rect 32116 26682 32172 26684
rect 32196 26682 32252 26684
rect 31956 26630 32002 26682
rect 32002 26630 32012 26682
rect 32036 26630 32066 26682
rect 32066 26630 32078 26682
rect 32078 26630 32092 26682
rect 32116 26630 32130 26682
rect 32130 26630 32142 26682
rect 32142 26630 32172 26682
rect 32196 26630 32206 26682
rect 32206 26630 32252 26682
rect 31956 26628 32012 26630
rect 32036 26628 32092 26630
rect 32116 26628 32172 26630
rect 32196 26628 32252 26630
rect 36956 26682 37012 26684
rect 37036 26682 37092 26684
rect 37116 26682 37172 26684
rect 37196 26682 37252 26684
rect 36956 26630 37002 26682
rect 37002 26630 37012 26682
rect 37036 26630 37066 26682
rect 37066 26630 37078 26682
rect 37078 26630 37092 26682
rect 37116 26630 37130 26682
rect 37130 26630 37142 26682
rect 37142 26630 37172 26682
rect 37196 26630 37206 26682
rect 37206 26630 37252 26682
rect 36956 26628 37012 26630
rect 37036 26628 37092 26630
rect 37116 26628 37172 26630
rect 37196 26628 37252 26630
rect 2616 26138 2672 26140
rect 2696 26138 2752 26140
rect 2776 26138 2832 26140
rect 2856 26138 2912 26140
rect 2616 26086 2662 26138
rect 2662 26086 2672 26138
rect 2696 26086 2726 26138
rect 2726 26086 2738 26138
rect 2738 26086 2752 26138
rect 2776 26086 2790 26138
rect 2790 26086 2802 26138
rect 2802 26086 2832 26138
rect 2856 26086 2866 26138
rect 2866 26086 2912 26138
rect 2616 26084 2672 26086
rect 2696 26084 2752 26086
rect 2776 26084 2832 26086
rect 2856 26084 2912 26086
rect 7616 26138 7672 26140
rect 7696 26138 7752 26140
rect 7776 26138 7832 26140
rect 7856 26138 7912 26140
rect 7616 26086 7662 26138
rect 7662 26086 7672 26138
rect 7696 26086 7726 26138
rect 7726 26086 7738 26138
rect 7738 26086 7752 26138
rect 7776 26086 7790 26138
rect 7790 26086 7802 26138
rect 7802 26086 7832 26138
rect 7856 26086 7866 26138
rect 7866 26086 7912 26138
rect 7616 26084 7672 26086
rect 7696 26084 7752 26086
rect 7776 26084 7832 26086
rect 7856 26084 7912 26086
rect 12616 26138 12672 26140
rect 12696 26138 12752 26140
rect 12776 26138 12832 26140
rect 12856 26138 12912 26140
rect 12616 26086 12662 26138
rect 12662 26086 12672 26138
rect 12696 26086 12726 26138
rect 12726 26086 12738 26138
rect 12738 26086 12752 26138
rect 12776 26086 12790 26138
rect 12790 26086 12802 26138
rect 12802 26086 12832 26138
rect 12856 26086 12866 26138
rect 12866 26086 12912 26138
rect 12616 26084 12672 26086
rect 12696 26084 12752 26086
rect 12776 26084 12832 26086
rect 12856 26084 12912 26086
rect 17616 26138 17672 26140
rect 17696 26138 17752 26140
rect 17776 26138 17832 26140
rect 17856 26138 17912 26140
rect 17616 26086 17662 26138
rect 17662 26086 17672 26138
rect 17696 26086 17726 26138
rect 17726 26086 17738 26138
rect 17738 26086 17752 26138
rect 17776 26086 17790 26138
rect 17790 26086 17802 26138
rect 17802 26086 17832 26138
rect 17856 26086 17866 26138
rect 17866 26086 17912 26138
rect 17616 26084 17672 26086
rect 17696 26084 17752 26086
rect 17776 26084 17832 26086
rect 17856 26084 17912 26086
rect 22616 26138 22672 26140
rect 22696 26138 22752 26140
rect 22776 26138 22832 26140
rect 22856 26138 22912 26140
rect 22616 26086 22662 26138
rect 22662 26086 22672 26138
rect 22696 26086 22726 26138
rect 22726 26086 22738 26138
rect 22738 26086 22752 26138
rect 22776 26086 22790 26138
rect 22790 26086 22802 26138
rect 22802 26086 22832 26138
rect 22856 26086 22866 26138
rect 22866 26086 22912 26138
rect 22616 26084 22672 26086
rect 22696 26084 22752 26086
rect 22776 26084 22832 26086
rect 22856 26084 22912 26086
rect 27616 26138 27672 26140
rect 27696 26138 27752 26140
rect 27776 26138 27832 26140
rect 27856 26138 27912 26140
rect 27616 26086 27662 26138
rect 27662 26086 27672 26138
rect 27696 26086 27726 26138
rect 27726 26086 27738 26138
rect 27738 26086 27752 26138
rect 27776 26086 27790 26138
rect 27790 26086 27802 26138
rect 27802 26086 27832 26138
rect 27856 26086 27866 26138
rect 27866 26086 27912 26138
rect 27616 26084 27672 26086
rect 27696 26084 27752 26086
rect 27776 26084 27832 26086
rect 27856 26084 27912 26086
rect 32616 26138 32672 26140
rect 32696 26138 32752 26140
rect 32776 26138 32832 26140
rect 32856 26138 32912 26140
rect 32616 26086 32662 26138
rect 32662 26086 32672 26138
rect 32696 26086 32726 26138
rect 32726 26086 32738 26138
rect 32738 26086 32752 26138
rect 32776 26086 32790 26138
rect 32790 26086 32802 26138
rect 32802 26086 32832 26138
rect 32856 26086 32866 26138
rect 32866 26086 32912 26138
rect 32616 26084 32672 26086
rect 32696 26084 32752 26086
rect 32776 26084 32832 26086
rect 32856 26084 32912 26086
rect 37616 26138 37672 26140
rect 37696 26138 37752 26140
rect 37776 26138 37832 26140
rect 37856 26138 37912 26140
rect 37616 26086 37662 26138
rect 37662 26086 37672 26138
rect 37696 26086 37726 26138
rect 37726 26086 37738 26138
rect 37738 26086 37752 26138
rect 37776 26086 37790 26138
rect 37790 26086 37802 26138
rect 37802 26086 37832 26138
rect 37856 26086 37866 26138
rect 37866 26086 37912 26138
rect 37616 26084 37672 26086
rect 37696 26084 37752 26086
rect 37776 26084 37832 26086
rect 37856 26084 37912 26086
rect 1956 25594 2012 25596
rect 2036 25594 2092 25596
rect 2116 25594 2172 25596
rect 2196 25594 2252 25596
rect 1956 25542 2002 25594
rect 2002 25542 2012 25594
rect 2036 25542 2066 25594
rect 2066 25542 2078 25594
rect 2078 25542 2092 25594
rect 2116 25542 2130 25594
rect 2130 25542 2142 25594
rect 2142 25542 2172 25594
rect 2196 25542 2206 25594
rect 2206 25542 2252 25594
rect 1956 25540 2012 25542
rect 2036 25540 2092 25542
rect 2116 25540 2172 25542
rect 2196 25540 2252 25542
rect 6956 25594 7012 25596
rect 7036 25594 7092 25596
rect 7116 25594 7172 25596
rect 7196 25594 7252 25596
rect 6956 25542 7002 25594
rect 7002 25542 7012 25594
rect 7036 25542 7066 25594
rect 7066 25542 7078 25594
rect 7078 25542 7092 25594
rect 7116 25542 7130 25594
rect 7130 25542 7142 25594
rect 7142 25542 7172 25594
rect 7196 25542 7206 25594
rect 7206 25542 7252 25594
rect 6956 25540 7012 25542
rect 7036 25540 7092 25542
rect 7116 25540 7172 25542
rect 7196 25540 7252 25542
rect 11956 25594 12012 25596
rect 12036 25594 12092 25596
rect 12116 25594 12172 25596
rect 12196 25594 12252 25596
rect 11956 25542 12002 25594
rect 12002 25542 12012 25594
rect 12036 25542 12066 25594
rect 12066 25542 12078 25594
rect 12078 25542 12092 25594
rect 12116 25542 12130 25594
rect 12130 25542 12142 25594
rect 12142 25542 12172 25594
rect 12196 25542 12206 25594
rect 12206 25542 12252 25594
rect 11956 25540 12012 25542
rect 12036 25540 12092 25542
rect 12116 25540 12172 25542
rect 12196 25540 12252 25542
rect 16956 25594 17012 25596
rect 17036 25594 17092 25596
rect 17116 25594 17172 25596
rect 17196 25594 17252 25596
rect 16956 25542 17002 25594
rect 17002 25542 17012 25594
rect 17036 25542 17066 25594
rect 17066 25542 17078 25594
rect 17078 25542 17092 25594
rect 17116 25542 17130 25594
rect 17130 25542 17142 25594
rect 17142 25542 17172 25594
rect 17196 25542 17206 25594
rect 17206 25542 17252 25594
rect 16956 25540 17012 25542
rect 17036 25540 17092 25542
rect 17116 25540 17172 25542
rect 17196 25540 17252 25542
rect 21956 25594 22012 25596
rect 22036 25594 22092 25596
rect 22116 25594 22172 25596
rect 22196 25594 22252 25596
rect 21956 25542 22002 25594
rect 22002 25542 22012 25594
rect 22036 25542 22066 25594
rect 22066 25542 22078 25594
rect 22078 25542 22092 25594
rect 22116 25542 22130 25594
rect 22130 25542 22142 25594
rect 22142 25542 22172 25594
rect 22196 25542 22206 25594
rect 22206 25542 22252 25594
rect 21956 25540 22012 25542
rect 22036 25540 22092 25542
rect 22116 25540 22172 25542
rect 22196 25540 22252 25542
rect 26956 25594 27012 25596
rect 27036 25594 27092 25596
rect 27116 25594 27172 25596
rect 27196 25594 27252 25596
rect 26956 25542 27002 25594
rect 27002 25542 27012 25594
rect 27036 25542 27066 25594
rect 27066 25542 27078 25594
rect 27078 25542 27092 25594
rect 27116 25542 27130 25594
rect 27130 25542 27142 25594
rect 27142 25542 27172 25594
rect 27196 25542 27206 25594
rect 27206 25542 27252 25594
rect 26956 25540 27012 25542
rect 27036 25540 27092 25542
rect 27116 25540 27172 25542
rect 27196 25540 27252 25542
rect 31956 25594 32012 25596
rect 32036 25594 32092 25596
rect 32116 25594 32172 25596
rect 32196 25594 32252 25596
rect 31956 25542 32002 25594
rect 32002 25542 32012 25594
rect 32036 25542 32066 25594
rect 32066 25542 32078 25594
rect 32078 25542 32092 25594
rect 32116 25542 32130 25594
rect 32130 25542 32142 25594
rect 32142 25542 32172 25594
rect 32196 25542 32206 25594
rect 32206 25542 32252 25594
rect 31956 25540 32012 25542
rect 32036 25540 32092 25542
rect 32116 25540 32172 25542
rect 32196 25540 32252 25542
rect 36956 25594 37012 25596
rect 37036 25594 37092 25596
rect 37116 25594 37172 25596
rect 37196 25594 37252 25596
rect 36956 25542 37002 25594
rect 37002 25542 37012 25594
rect 37036 25542 37066 25594
rect 37066 25542 37078 25594
rect 37078 25542 37092 25594
rect 37116 25542 37130 25594
rect 37130 25542 37142 25594
rect 37142 25542 37172 25594
rect 37196 25542 37206 25594
rect 37206 25542 37252 25594
rect 36956 25540 37012 25542
rect 37036 25540 37092 25542
rect 37116 25540 37172 25542
rect 37196 25540 37252 25542
rect 2616 25050 2672 25052
rect 2696 25050 2752 25052
rect 2776 25050 2832 25052
rect 2856 25050 2912 25052
rect 2616 24998 2662 25050
rect 2662 24998 2672 25050
rect 2696 24998 2726 25050
rect 2726 24998 2738 25050
rect 2738 24998 2752 25050
rect 2776 24998 2790 25050
rect 2790 24998 2802 25050
rect 2802 24998 2832 25050
rect 2856 24998 2866 25050
rect 2866 24998 2912 25050
rect 2616 24996 2672 24998
rect 2696 24996 2752 24998
rect 2776 24996 2832 24998
rect 2856 24996 2912 24998
rect 7616 25050 7672 25052
rect 7696 25050 7752 25052
rect 7776 25050 7832 25052
rect 7856 25050 7912 25052
rect 7616 24998 7662 25050
rect 7662 24998 7672 25050
rect 7696 24998 7726 25050
rect 7726 24998 7738 25050
rect 7738 24998 7752 25050
rect 7776 24998 7790 25050
rect 7790 24998 7802 25050
rect 7802 24998 7832 25050
rect 7856 24998 7866 25050
rect 7866 24998 7912 25050
rect 7616 24996 7672 24998
rect 7696 24996 7752 24998
rect 7776 24996 7832 24998
rect 7856 24996 7912 24998
rect 12616 25050 12672 25052
rect 12696 25050 12752 25052
rect 12776 25050 12832 25052
rect 12856 25050 12912 25052
rect 12616 24998 12662 25050
rect 12662 24998 12672 25050
rect 12696 24998 12726 25050
rect 12726 24998 12738 25050
rect 12738 24998 12752 25050
rect 12776 24998 12790 25050
rect 12790 24998 12802 25050
rect 12802 24998 12832 25050
rect 12856 24998 12866 25050
rect 12866 24998 12912 25050
rect 12616 24996 12672 24998
rect 12696 24996 12752 24998
rect 12776 24996 12832 24998
rect 12856 24996 12912 24998
rect 17616 25050 17672 25052
rect 17696 25050 17752 25052
rect 17776 25050 17832 25052
rect 17856 25050 17912 25052
rect 17616 24998 17662 25050
rect 17662 24998 17672 25050
rect 17696 24998 17726 25050
rect 17726 24998 17738 25050
rect 17738 24998 17752 25050
rect 17776 24998 17790 25050
rect 17790 24998 17802 25050
rect 17802 24998 17832 25050
rect 17856 24998 17866 25050
rect 17866 24998 17912 25050
rect 17616 24996 17672 24998
rect 17696 24996 17752 24998
rect 17776 24996 17832 24998
rect 17856 24996 17912 24998
rect 22616 25050 22672 25052
rect 22696 25050 22752 25052
rect 22776 25050 22832 25052
rect 22856 25050 22912 25052
rect 22616 24998 22662 25050
rect 22662 24998 22672 25050
rect 22696 24998 22726 25050
rect 22726 24998 22738 25050
rect 22738 24998 22752 25050
rect 22776 24998 22790 25050
rect 22790 24998 22802 25050
rect 22802 24998 22832 25050
rect 22856 24998 22866 25050
rect 22866 24998 22912 25050
rect 22616 24996 22672 24998
rect 22696 24996 22752 24998
rect 22776 24996 22832 24998
rect 22856 24996 22912 24998
rect 27616 25050 27672 25052
rect 27696 25050 27752 25052
rect 27776 25050 27832 25052
rect 27856 25050 27912 25052
rect 27616 24998 27662 25050
rect 27662 24998 27672 25050
rect 27696 24998 27726 25050
rect 27726 24998 27738 25050
rect 27738 24998 27752 25050
rect 27776 24998 27790 25050
rect 27790 24998 27802 25050
rect 27802 24998 27832 25050
rect 27856 24998 27866 25050
rect 27866 24998 27912 25050
rect 27616 24996 27672 24998
rect 27696 24996 27752 24998
rect 27776 24996 27832 24998
rect 27856 24996 27912 24998
rect 32616 25050 32672 25052
rect 32696 25050 32752 25052
rect 32776 25050 32832 25052
rect 32856 25050 32912 25052
rect 32616 24998 32662 25050
rect 32662 24998 32672 25050
rect 32696 24998 32726 25050
rect 32726 24998 32738 25050
rect 32738 24998 32752 25050
rect 32776 24998 32790 25050
rect 32790 24998 32802 25050
rect 32802 24998 32832 25050
rect 32856 24998 32866 25050
rect 32866 24998 32912 25050
rect 32616 24996 32672 24998
rect 32696 24996 32752 24998
rect 32776 24996 32832 24998
rect 32856 24996 32912 24998
rect 37616 25050 37672 25052
rect 37696 25050 37752 25052
rect 37776 25050 37832 25052
rect 37856 25050 37912 25052
rect 37616 24998 37662 25050
rect 37662 24998 37672 25050
rect 37696 24998 37726 25050
rect 37726 24998 37738 25050
rect 37738 24998 37752 25050
rect 37776 24998 37790 25050
rect 37790 24998 37802 25050
rect 37802 24998 37832 25050
rect 37856 24998 37866 25050
rect 37866 24998 37912 25050
rect 37616 24996 37672 24998
rect 37696 24996 37752 24998
rect 37776 24996 37832 24998
rect 37856 24996 37912 24998
rect 1956 24506 2012 24508
rect 2036 24506 2092 24508
rect 2116 24506 2172 24508
rect 2196 24506 2252 24508
rect 1956 24454 2002 24506
rect 2002 24454 2012 24506
rect 2036 24454 2066 24506
rect 2066 24454 2078 24506
rect 2078 24454 2092 24506
rect 2116 24454 2130 24506
rect 2130 24454 2142 24506
rect 2142 24454 2172 24506
rect 2196 24454 2206 24506
rect 2206 24454 2252 24506
rect 1956 24452 2012 24454
rect 2036 24452 2092 24454
rect 2116 24452 2172 24454
rect 2196 24452 2252 24454
rect 6956 24506 7012 24508
rect 7036 24506 7092 24508
rect 7116 24506 7172 24508
rect 7196 24506 7252 24508
rect 6956 24454 7002 24506
rect 7002 24454 7012 24506
rect 7036 24454 7066 24506
rect 7066 24454 7078 24506
rect 7078 24454 7092 24506
rect 7116 24454 7130 24506
rect 7130 24454 7142 24506
rect 7142 24454 7172 24506
rect 7196 24454 7206 24506
rect 7206 24454 7252 24506
rect 6956 24452 7012 24454
rect 7036 24452 7092 24454
rect 7116 24452 7172 24454
rect 7196 24452 7252 24454
rect 11956 24506 12012 24508
rect 12036 24506 12092 24508
rect 12116 24506 12172 24508
rect 12196 24506 12252 24508
rect 11956 24454 12002 24506
rect 12002 24454 12012 24506
rect 12036 24454 12066 24506
rect 12066 24454 12078 24506
rect 12078 24454 12092 24506
rect 12116 24454 12130 24506
rect 12130 24454 12142 24506
rect 12142 24454 12172 24506
rect 12196 24454 12206 24506
rect 12206 24454 12252 24506
rect 11956 24452 12012 24454
rect 12036 24452 12092 24454
rect 12116 24452 12172 24454
rect 12196 24452 12252 24454
rect 16956 24506 17012 24508
rect 17036 24506 17092 24508
rect 17116 24506 17172 24508
rect 17196 24506 17252 24508
rect 16956 24454 17002 24506
rect 17002 24454 17012 24506
rect 17036 24454 17066 24506
rect 17066 24454 17078 24506
rect 17078 24454 17092 24506
rect 17116 24454 17130 24506
rect 17130 24454 17142 24506
rect 17142 24454 17172 24506
rect 17196 24454 17206 24506
rect 17206 24454 17252 24506
rect 16956 24452 17012 24454
rect 17036 24452 17092 24454
rect 17116 24452 17172 24454
rect 17196 24452 17252 24454
rect 21956 24506 22012 24508
rect 22036 24506 22092 24508
rect 22116 24506 22172 24508
rect 22196 24506 22252 24508
rect 21956 24454 22002 24506
rect 22002 24454 22012 24506
rect 22036 24454 22066 24506
rect 22066 24454 22078 24506
rect 22078 24454 22092 24506
rect 22116 24454 22130 24506
rect 22130 24454 22142 24506
rect 22142 24454 22172 24506
rect 22196 24454 22206 24506
rect 22206 24454 22252 24506
rect 21956 24452 22012 24454
rect 22036 24452 22092 24454
rect 22116 24452 22172 24454
rect 22196 24452 22252 24454
rect 26956 24506 27012 24508
rect 27036 24506 27092 24508
rect 27116 24506 27172 24508
rect 27196 24506 27252 24508
rect 26956 24454 27002 24506
rect 27002 24454 27012 24506
rect 27036 24454 27066 24506
rect 27066 24454 27078 24506
rect 27078 24454 27092 24506
rect 27116 24454 27130 24506
rect 27130 24454 27142 24506
rect 27142 24454 27172 24506
rect 27196 24454 27206 24506
rect 27206 24454 27252 24506
rect 26956 24452 27012 24454
rect 27036 24452 27092 24454
rect 27116 24452 27172 24454
rect 27196 24452 27252 24454
rect 31956 24506 32012 24508
rect 32036 24506 32092 24508
rect 32116 24506 32172 24508
rect 32196 24506 32252 24508
rect 31956 24454 32002 24506
rect 32002 24454 32012 24506
rect 32036 24454 32066 24506
rect 32066 24454 32078 24506
rect 32078 24454 32092 24506
rect 32116 24454 32130 24506
rect 32130 24454 32142 24506
rect 32142 24454 32172 24506
rect 32196 24454 32206 24506
rect 32206 24454 32252 24506
rect 31956 24452 32012 24454
rect 32036 24452 32092 24454
rect 32116 24452 32172 24454
rect 32196 24452 32252 24454
rect 36956 24506 37012 24508
rect 37036 24506 37092 24508
rect 37116 24506 37172 24508
rect 37196 24506 37252 24508
rect 36956 24454 37002 24506
rect 37002 24454 37012 24506
rect 37036 24454 37066 24506
rect 37066 24454 37078 24506
rect 37078 24454 37092 24506
rect 37116 24454 37130 24506
rect 37130 24454 37142 24506
rect 37142 24454 37172 24506
rect 37196 24454 37206 24506
rect 37206 24454 37252 24506
rect 36956 24452 37012 24454
rect 37036 24452 37092 24454
rect 37116 24452 37172 24454
rect 37196 24452 37252 24454
rect 2616 23962 2672 23964
rect 2696 23962 2752 23964
rect 2776 23962 2832 23964
rect 2856 23962 2912 23964
rect 2616 23910 2662 23962
rect 2662 23910 2672 23962
rect 2696 23910 2726 23962
rect 2726 23910 2738 23962
rect 2738 23910 2752 23962
rect 2776 23910 2790 23962
rect 2790 23910 2802 23962
rect 2802 23910 2832 23962
rect 2856 23910 2866 23962
rect 2866 23910 2912 23962
rect 2616 23908 2672 23910
rect 2696 23908 2752 23910
rect 2776 23908 2832 23910
rect 2856 23908 2912 23910
rect 7616 23962 7672 23964
rect 7696 23962 7752 23964
rect 7776 23962 7832 23964
rect 7856 23962 7912 23964
rect 7616 23910 7662 23962
rect 7662 23910 7672 23962
rect 7696 23910 7726 23962
rect 7726 23910 7738 23962
rect 7738 23910 7752 23962
rect 7776 23910 7790 23962
rect 7790 23910 7802 23962
rect 7802 23910 7832 23962
rect 7856 23910 7866 23962
rect 7866 23910 7912 23962
rect 7616 23908 7672 23910
rect 7696 23908 7752 23910
rect 7776 23908 7832 23910
rect 7856 23908 7912 23910
rect 12616 23962 12672 23964
rect 12696 23962 12752 23964
rect 12776 23962 12832 23964
rect 12856 23962 12912 23964
rect 12616 23910 12662 23962
rect 12662 23910 12672 23962
rect 12696 23910 12726 23962
rect 12726 23910 12738 23962
rect 12738 23910 12752 23962
rect 12776 23910 12790 23962
rect 12790 23910 12802 23962
rect 12802 23910 12832 23962
rect 12856 23910 12866 23962
rect 12866 23910 12912 23962
rect 12616 23908 12672 23910
rect 12696 23908 12752 23910
rect 12776 23908 12832 23910
rect 12856 23908 12912 23910
rect 17616 23962 17672 23964
rect 17696 23962 17752 23964
rect 17776 23962 17832 23964
rect 17856 23962 17912 23964
rect 17616 23910 17662 23962
rect 17662 23910 17672 23962
rect 17696 23910 17726 23962
rect 17726 23910 17738 23962
rect 17738 23910 17752 23962
rect 17776 23910 17790 23962
rect 17790 23910 17802 23962
rect 17802 23910 17832 23962
rect 17856 23910 17866 23962
rect 17866 23910 17912 23962
rect 17616 23908 17672 23910
rect 17696 23908 17752 23910
rect 17776 23908 17832 23910
rect 17856 23908 17912 23910
rect 22616 23962 22672 23964
rect 22696 23962 22752 23964
rect 22776 23962 22832 23964
rect 22856 23962 22912 23964
rect 22616 23910 22662 23962
rect 22662 23910 22672 23962
rect 22696 23910 22726 23962
rect 22726 23910 22738 23962
rect 22738 23910 22752 23962
rect 22776 23910 22790 23962
rect 22790 23910 22802 23962
rect 22802 23910 22832 23962
rect 22856 23910 22866 23962
rect 22866 23910 22912 23962
rect 22616 23908 22672 23910
rect 22696 23908 22752 23910
rect 22776 23908 22832 23910
rect 22856 23908 22912 23910
rect 27616 23962 27672 23964
rect 27696 23962 27752 23964
rect 27776 23962 27832 23964
rect 27856 23962 27912 23964
rect 27616 23910 27662 23962
rect 27662 23910 27672 23962
rect 27696 23910 27726 23962
rect 27726 23910 27738 23962
rect 27738 23910 27752 23962
rect 27776 23910 27790 23962
rect 27790 23910 27802 23962
rect 27802 23910 27832 23962
rect 27856 23910 27866 23962
rect 27866 23910 27912 23962
rect 27616 23908 27672 23910
rect 27696 23908 27752 23910
rect 27776 23908 27832 23910
rect 27856 23908 27912 23910
rect 32616 23962 32672 23964
rect 32696 23962 32752 23964
rect 32776 23962 32832 23964
rect 32856 23962 32912 23964
rect 32616 23910 32662 23962
rect 32662 23910 32672 23962
rect 32696 23910 32726 23962
rect 32726 23910 32738 23962
rect 32738 23910 32752 23962
rect 32776 23910 32790 23962
rect 32790 23910 32802 23962
rect 32802 23910 32832 23962
rect 32856 23910 32866 23962
rect 32866 23910 32912 23962
rect 32616 23908 32672 23910
rect 32696 23908 32752 23910
rect 32776 23908 32832 23910
rect 32856 23908 32912 23910
rect 37616 23962 37672 23964
rect 37696 23962 37752 23964
rect 37776 23962 37832 23964
rect 37856 23962 37912 23964
rect 37616 23910 37662 23962
rect 37662 23910 37672 23962
rect 37696 23910 37726 23962
rect 37726 23910 37738 23962
rect 37738 23910 37752 23962
rect 37776 23910 37790 23962
rect 37790 23910 37802 23962
rect 37802 23910 37832 23962
rect 37856 23910 37866 23962
rect 37866 23910 37912 23962
rect 37616 23908 37672 23910
rect 37696 23908 37752 23910
rect 37776 23908 37832 23910
rect 37856 23908 37912 23910
rect 1956 23418 2012 23420
rect 2036 23418 2092 23420
rect 2116 23418 2172 23420
rect 2196 23418 2252 23420
rect 1956 23366 2002 23418
rect 2002 23366 2012 23418
rect 2036 23366 2066 23418
rect 2066 23366 2078 23418
rect 2078 23366 2092 23418
rect 2116 23366 2130 23418
rect 2130 23366 2142 23418
rect 2142 23366 2172 23418
rect 2196 23366 2206 23418
rect 2206 23366 2252 23418
rect 1956 23364 2012 23366
rect 2036 23364 2092 23366
rect 2116 23364 2172 23366
rect 2196 23364 2252 23366
rect 6956 23418 7012 23420
rect 7036 23418 7092 23420
rect 7116 23418 7172 23420
rect 7196 23418 7252 23420
rect 6956 23366 7002 23418
rect 7002 23366 7012 23418
rect 7036 23366 7066 23418
rect 7066 23366 7078 23418
rect 7078 23366 7092 23418
rect 7116 23366 7130 23418
rect 7130 23366 7142 23418
rect 7142 23366 7172 23418
rect 7196 23366 7206 23418
rect 7206 23366 7252 23418
rect 6956 23364 7012 23366
rect 7036 23364 7092 23366
rect 7116 23364 7172 23366
rect 7196 23364 7252 23366
rect 11956 23418 12012 23420
rect 12036 23418 12092 23420
rect 12116 23418 12172 23420
rect 12196 23418 12252 23420
rect 11956 23366 12002 23418
rect 12002 23366 12012 23418
rect 12036 23366 12066 23418
rect 12066 23366 12078 23418
rect 12078 23366 12092 23418
rect 12116 23366 12130 23418
rect 12130 23366 12142 23418
rect 12142 23366 12172 23418
rect 12196 23366 12206 23418
rect 12206 23366 12252 23418
rect 11956 23364 12012 23366
rect 12036 23364 12092 23366
rect 12116 23364 12172 23366
rect 12196 23364 12252 23366
rect 16956 23418 17012 23420
rect 17036 23418 17092 23420
rect 17116 23418 17172 23420
rect 17196 23418 17252 23420
rect 16956 23366 17002 23418
rect 17002 23366 17012 23418
rect 17036 23366 17066 23418
rect 17066 23366 17078 23418
rect 17078 23366 17092 23418
rect 17116 23366 17130 23418
rect 17130 23366 17142 23418
rect 17142 23366 17172 23418
rect 17196 23366 17206 23418
rect 17206 23366 17252 23418
rect 16956 23364 17012 23366
rect 17036 23364 17092 23366
rect 17116 23364 17172 23366
rect 17196 23364 17252 23366
rect 21956 23418 22012 23420
rect 22036 23418 22092 23420
rect 22116 23418 22172 23420
rect 22196 23418 22252 23420
rect 21956 23366 22002 23418
rect 22002 23366 22012 23418
rect 22036 23366 22066 23418
rect 22066 23366 22078 23418
rect 22078 23366 22092 23418
rect 22116 23366 22130 23418
rect 22130 23366 22142 23418
rect 22142 23366 22172 23418
rect 22196 23366 22206 23418
rect 22206 23366 22252 23418
rect 21956 23364 22012 23366
rect 22036 23364 22092 23366
rect 22116 23364 22172 23366
rect 22196 23364 22252 23366
rect 26956 23418 27012 23420
rect 27036 23418 27092 23420
rect 27116 23418 27172 23420
rect 27196 23418 27252 23420
rect 26956 23366 27002 23418
rect 27002 23366 27012 23418
rect 27036 23366 27066 23418
rect 27066 23366 27078 23418
rect 27078 23366 27092 23418
rect 27116 23366 27130 23418
rect 27130 23366 27142 23418
rect 27142 23366 27172 23418
rect 27196 23366 27206 23418
rect 27206 23366 27252 23418
rect 26956 23364 27012 23366
rect 27036 23364 27092 23366
rect 27116 23364 27172 23366
rect 27196 23364 27252 23366
rect 31956 23418 32012 23420
rect 32036 23418 32092 23420
rect 32116 23418 32172 23420
rect 32196 23418 32252 23420
rect 31956 23366 32002 23418
rect 32002 23366 32012 23418
rect 32036 23366 32066 23418
rect 32066 23366 32078 23418
rect 32078 23366 32092 23418
rect 32116 23366 32130 23418
rect 32130 23366 32142 23418
rect 32142 23366 32172 23418
rect 32196 23366 32206 23418
rect 32206 23366 32252 23418
rect 31956 23364 32012 23366
rect 32036 23364 32092 23366
rect 32116 23364 32172 23366
rect 32196 23364 32252 23366
rect 36956 23418 37012 23420
rect 37036 23418 37092 23420
rect 37116 23418 37172 23420
rect 37196 23418 37252 23420
rect 36956 23366 37002 23418
rect 37002 23366 37012 23418
rect 37036 23366 37066 23418
rect 37066 23366 37078 23418
rect 37078 23366 37092 23418
rect 37116 23366 37130 23418
rect 37130 23366 37142 23418
rect 37142 23366 37172 23418
rect 37196 23366 37206 23418
rect 37206 23366 37252 23418
rect 36956 23364 37012 23366
rect 37036 23364 37092 23366
rect 37116 23364 37172 23366
rect 37196 23364 37252 23366
rect 2616 22874 2672 22876
rect 2696 22874 2752 22876
rect 2776 22874 2832 22876
rect 2856 22874 2912 22876
rect 2616 22822 2662 22874
rect 2662 22822 2672 22874
rect 2696 22822 2726 22874
rect 2726 22822 2738 22874
rect 2738 22822 2752 22874
rect 2776 22822 2790 22874
rect 2790 22822 2802 22874
rect 2802 22822 2832 22874
rect 2856 22822 2866 22874
rect 2866 22822 2912 22874
rect 2616 22820 2672 22822
rect 2696 22820 2752 22822
rect 2776 22820 2832 22822
rect 2856 22820 2912 22822
rect 7616 22874 7672 22876
rect 7696 22874 7752 22876
rect 7776 22874 7832 22876
rect 7856 22874 7912 22876
rect 7616 22822 7662 22874
rect 7662 22822 7672 22874
rect 7696 22822 7726 22874
rect 7726 22822 7738 22874
rect 7738 22822 7752 22874
rect 7776 22822 7790 22874
rect 7790 22822 7802 22874
rect 7802 22822 7832 22874
rect 7856 22822 7866 22874
rect 7866 22822 7912 22874
rect 7616 22820 7672 22822
rect 7696 22820 7752 22822
rect 7776 22820 7832 22822
rect 7856 22820 7912 22822
rect 12616 22874 12672 22876
rect 12696 22874 12752 22876
rect 12776 22874 12832 22876
rect 12856 22874 12912 22876
rect 12616 22822 12662 22874
rect 12662 22822 12672 22874
rect 12696 22822 12726 22874
rect 12726 22822 12738 22874
rect 12738 22822 12752 22874
rect 12776 22822 12790 22874
rect 12790 22822 12802 22874
rect 12802 22822 12832 22874
rect 12856 22822 12866 22874
rect 12866 22822 12912 22874
rect 12616 22820 12672 22822
rect 12696 22820 12752 22822
rect 12776 22820 12832 22822
rect 12856 22820 12912 22822
rect 17616 22874 17672 22876
rect 17696 22874 17752 22876
rect 17776 22874 17832 22876
rect 17856 22874 17912 22876
rect 17616 22822 17662 22874
rect 17662 22822 17672 22874
rect 17696 22822 17726 22874
rect 17726 22822 17738 22874
rect 17738 22822 17752 22874
rect 17776 22822 17790 22874
rect 17790 22822 17802 22874
rect 17802 22822 17832 22874
rect 17856 22822 17866 22874
rect 17866 22822 17912 22874
rect 17616 22820 17672 22822
rect 17696 22820 17752 22822
rect 17776 22820 17832 22822
rect 17856 22820 17912 22822
rect 22616 22874 22672 22876
rect 22696 22874 22752 22876
rect 22776 22874 22832 22876
rect 22856 22874 22912 22876
rect 22616 22822 22662 22874
rect 22662 22822 22672 22874
rect 22696 22822 22726 22874
rect 22726 22822 22738 22874
rect 22738 22822 22752 22874
rect 22776 22822 22790 22874
rect 22790 22822 22802 22874
rect 22802 22822 22832 22874
rect 22856 22822 22866 22874
rect 22866 22822 22912 22874
rect 22616 22820 22672 22822
rect 22696 22820 22752 22822
rect 22776 22820 22832 22822
rect 22856 22820 22912 22822
rect 27616 22874 27672 22876
rect 27696 22874 27752 22876
rect 27776 22874 27832 22876
rect 27856 22874 27912 22876
rect 27616 22822 27662 22874
rect 27662 22822 27672 22874
rect 27696 22822 27726 22874
rect 27726 22822 27738 22874
rect 27738 22822 27752 22874
rect 27776 22822 27790 22874
rect 27790 22822 27802 22874
rect 27802 22822 27832 22874
rect 27856 22822 27866 22874
rect 27866 22822 27912 22874
rect 27616 22820 27672 22822
rect 27696 22820 27752 22822
rect 27776 22820 27832 22822
rect 27856 22820 27912 22822
rect 32616 22874 32672 22876
rect 32696 22874 32752 22876
rect 32776 22874 32832 22876
rect 32856 22874 32912 22876
rect 32616 22822 32662 22874
rect 32662 22822 32672 22874
rect 32696 22822 32726 22874
rect 32726 22822 32738 22874
rect 32738 22822 32752 22874
rect 32776 22822 32790 22874
rect 32790 22822 32802 22874
rect 32802 22822 32832 22874
rect 32856 22822 32866 22874
rect 32866 22822 32912 22874
rect 32616 22820 32672 22822
rect 32696 22820 32752 22822
rect 32776 22820 32832 22822
rect 32856 22820 32912 22822
rect 37616 22874 37672 22876
rect 37696 22874 37752 22876
rect 37776 22874 37832 22876
rect 37856 22874 37912 22876
rect 37616 22822 37662 22874
rect 37662 22822 37672 22874
rect 37696 22822 37726 22874
rect 37726 22822 37738 22874
rect 37738 22822 37752 22874
rect 37776 22822 37790 22874
rect 37790 22822 37802 22874
rect 37802 22822 37832 22874
rect 37856 22822 37866 22874
rect 37866 22822 37912 22874
rect 37616 22820 37672 22822
rect 37696 22820 37752 22822
rect 37776 22820 37832 22822
rect 37856 22820 37912 22822
rect 1956 22330 2012 22332
rect 2036 22330 2092 22332
rect 2116 22330 2172 22332
rect 2196 22330 2252 22332
rect 1956 22278 2002 22330
rect 2002 22278 2012 22330
rect 2036 22278 2066 22330
rect 2066 22278 2078 22330
rect 2078 22278 2092 22330
rect 2116 22278 2130 22330
rect 2130 22278 2142 22330
rect 2142 22278 2172 22330
rect 2196 22278 2206 22330
rect 2206 22278 2252 22330
rect 1956 22276 2012 22278
rect 2036 22276 2092 22278
rect 2116 22276 2172 22278
rect 2196 22276 2252 22278
rect 6956 22330 7012 22332
rect 7036 22330 7092 22332
rect 7116 22330 7172 22332
rect 7196 22330 7252 22332
rect 6956 22278 7002 22330
rect 7002 22278 7012 22330
rect 7036 22278 7066 22330
rect 7066 22278 7078 22330
rect 7078 22278 7092 22330
rect 7116 22278 7130 22330
rect 7130 22278 7142 22330
rect 7142 22278 7172 22330
rect 7196 22278 7206 22330
rect 7206 22278 7252 22330
rect 6956 22276 7012 22278
rect 7036 22276 7092 22278
rect 7116 22276 7172 22278
rect 7196 22276 7252 22278
rect 11956 22330 12012 22332
rect 12036 22330 12092 22332
rect 12116 22330 12172 22332
rect 12196 22330 12252 22332
rect 11956 22278 12002 22330
rect 12002 22278 12012 22330
rect 12036 22278 12066 22330
rect 12066 22278 12078 22330
rect 12078 22278 12092 22330
rect 12116 22278 12130 22330
rect 12130 22278 12142 22330
rect 12142 22278 12172 22330
rect 12196 22278 12206 22330
rect 12206 22278 12252 22330
rect 11956 22276 12012 22278
rect 12036 22276 12092 22278
rect 12116 22276 12172 22278
rect 12196 22276 12252 22278
rect 16956 22330 17012 22332
rect 17036 22330 17092 22332
rect 17116 22330 17172 22332
rect 17196 22330 17252 22332
rect 16956 22278 17002 22330
rect 17002 22278 17012 22330
rect 17036 22278 17066 22330
rect 17066 22278 17078 22330
rect 17078 22278 17092 22330
rect 17116 22278 17130 22330
rect 17130 22278 17142 22330
rect 17142 22278 17172 22330
rect 17196 22278 17206 22330
rect 17206 22278 17252 22330
rect 16956 22276 17012 22278
rect 17036 22276 17092 22278
rect 17116 22276 17172 22278
rect 17196 22276 17252 22278
rect 21956 22330 22012 22332
rect 22036 22330 22092 22332
rect 22116 22330 22172 22332
rect 22196 22330 22252 22332
rect 21956 22278 22002 22330
rect 22002 22278 22012 22330
rect 22036 22278 22066 22330
rect 22066 22278 22078 22330
rect 22078 22278 22092 22330
rect 22116 22278 22130 22330
rect 22130 22278 22142 22330
rect 22142 22278 22172 22330
rect 22196 22278 22206 22330
rect 22206 22278 22252 22330
rect 21956 22276 22012 22278
rect 22036 22276 22092 22278
rect 22116 22276 22172 22278
rect 22196 22276 22252 22278
rect 26956 22330 27012 22332
rect 27036 22330 27092 22332
rect 27116 22330 27172 22332
rect 27196 22330 27252 22332
rect 26956 22278 27002 22330
rect 27002 22278 27012 22330
rect 27036 22278 27066 22330
rect 27066 22278 27078 22330
rect 27078 22278 27092 22330
rect 27116 22278 27130 22330
rect 27130 22278 27142 22330
rect 27142 22278 27172 22330
rect 27196 22278 27206 22330
rect 27206 22278 27252 22330
rect 26956 22276 27012 22278
rect 27036 22276 27092 22278
rect 27116 22276 27172 22278
rect 27196 22276 27252 22278
rect 31956 22330 32012 22332
rect 32036 22330 32092 22332
rect 32116 22330 32172 22332
rect 32196 22330 32252 22332
rect 31956 22278 32002 22330
rect 32002 22278 32012 22330
rect 32036 22278 32066 22330
rect 32066 22278 32078 22330
rect 32078 22278 32092 22330
rect 32116 22278 32130 22330
rect 32130 22278 32142 22330
rect 32142 22278 32172 22330
rect 32196 22278 32206 22330
rect 32206 22278 32252 22330
rect 31956 22276 32012 22278
rect 32036 22276 32092 22278
rect 32116 22276 32172 22278
rect 32196 22276 32252 22278
rect 36956 22330 37012 22332
rect 37036 22330 37092 22332
rect 37116 22330 37172 22332
rect 37196 22330 37252 22332
rect 36956 22278 37002 22330
rect 37002 22278 37012 22330
rect 37036 22278 37066 22330
rect 37066 22278 37078 22330
rect 37078 22278 37092 22330
rect 37116 22278 37130 22330
rect 37130 22278 37142 22330
rect 37142 22278 37172 22330
rect 37196 22278 37206 22330
rect 37206 22278 37252 22330
rect 36956 22276 37012 22278
rect 37036 22276 37092 22278
rect 37116 22276 37172 22278
rect 37196 22276 37252 22278
rect 2616 21786 2672 21788
rect 2696 21786 2752 21788
rect 2776 21786 2832 21788
rect 2856 21786 2912 21788
rect 2616 21734 2662 21786
rect 2662 21734 2672 21786
rect 2696 21734 2726 21786
rect 2726 21734 2738 21786
rect 2738 21734 2752 21786
rect 2776 21734 2790 21786
rect 2790 21734 2802 21786
rect 2802 21734 2832 21786
rect 2856 21734 2866 21786
rect 2866 21734 2912 21786
rect 2616 21732 2672 21734
rect 2696 21732 2752 21734
rect 2776 21732 2832 21734
rect 2856 21732 2912 21734
rect 7616 21786 7672 21788
rect 7696 21786 7752 21788
rect 7776 21786 7832 21788
rect 7856 21786 7912 21788
rect 7616 21734 7662 21786
rect 7662 21734 7672 21786
rect 7696 21734 7726 21786
rect 7726 21734 7738 21786
rect 7738 21734 7752 21786
rect 7776 21734 7790 21786
rect 7790 21734 7802 21786
rect 7802 21734 7832 21786
rect 7856 21734 7866 21786
rect 7866 21734 7912 21786
rect 7616 21732 7672 21734
rect 7696 21732 7752 21734
rect 7776 21732 7832 21734
rect 7856 21732 7912 21734
rect 12616 21786 12672 21788
rect 12696 21786 12752 21788
rect 12776 21786 12832 21788
rect 12856 21786 12912 21788
rect 12616 21734 12662 21786
rect 12662 21734 12672 21786
rect 12696 21734 12726 21786
rect 12726 21734 12738 21786
rect 12738 21734 12752 21786
rect 12776 21734 12790 21786
rect 12790 21734 12802 21786
rect 12802 21734 12832 21786
rect 12856 21734 12866 21786
rect 12866 21734 12912 21786
rect 12616 21732 12672 21734
rect 12696 21732 12752 21734
rect 12776 21732 12832 21734
rect 12856 21732 12912 21734
rect 17616 21786 17672 21788
rect 17696 21786 17752 21788
rect 17776 21786 17832 21788
rect 17856 21786 17912 21788
rect 17616 21734 17662 21786
rect 17662 21734 17672 21786
rect 17696 21734 17726 21786
rect 17726 21734 17738 21786
rect 17738 21734 17752 21786
rect 17776 21734 17790 21786
rect 17790 21734 17802 21786
rect 17802 21734 17832 21786
rect 17856 21734 17866 21786
rect 17866 21734 17912 21786
rect 17616 21732 17672 21734
rect 17696 21732 17752 21734
rect 17776 21732 17832 21734
rect 17856 21732 17912 21734
rect 22616 21786 22672 21788
rect 22696 21786 22752 21788
rect 22776 21786 22832 21788
rect 22856 21786 22912 21788
rect 22616 21734 22662 21786
rect 22662 21734 22672 21786
rect 22696 21734 22726 21786
rect 22726 21734 22738 21786
rect 22738 21734 22752 21786
rect 22776 21734 22790 21786
rect 22790 21734 22802 21786
rect 22802 21734 22832 21786
rect 22856 21734 22866 21786
rect 22866 21734 22912 21786
rect 22616 21732 22672 21734
rect 22696 21732 22752 21734
rect 22776 21732 22832 21734
rect 22856 21732 22912 21734
rect 27616 21786 27672 21788
rect 27696 21786 27752 21788
rect 27776 21786 27832 21788
rect 27856 21786 27912 21788
rect 27616 21734 27662 21786
rect 27662 21734 27672 21786
rect 27696 21734 27726 21786
rect 27726 21734 27738 21786
rect 27738 21734 27752 21786
rect 27776 21734 27790 21786
rect 27790 21734 27802 21786
rect 27802 21734 27832 21786
rect 27856 21734 27866 21786
rect 27866 21734 27912 21786
rect 27616 21732 27672 21734
rect 27696 21732 27752 21734
rect 27776 21732 27832 21734
rect 27856 21732 27912 21734
rect 32616 21786 32672 21788
rect 32696 21786 32752 21788
rect 32776 21786 32832 21788
rect 32856 21786 32912 21788
rect 32616 21734 32662 21786
rect 32662 21734 32672 21786
rect 32696 21734 32726 21786
rect 32726 21734 32738 21786
rect 32738 21734 32752 21786
rect 32776 21734 32790 21786
rect 32790 21734 32802 21786
rect 32802 21734 32832 21786
rect 32856 21734 32866 21786
rect 32866 21734 32912 21786
rect 32616 21732 32672 21734
rect 32696 21732 32752 21734
rect 32776 21732 32832 21734
rect 32856 21732 32912 21734
rect 938 21120 994 21176
rect 1956 21242 2012 21244
rect 2036 21242 2092 21244
rect 2116 21242 2172 21244
rect 2196 21242 2252 21244
rect 1956 21190 2002 21242
rect 2002 21190 2012 21242
rect 2036 21190 2066 21242
rect 2066 21190 2078 21242
rect 2078 21190 2092 21242
rect 2116 21190 2130 21242
rect 2130 21190 2142 21242
rect 2142 21190 2172 21242
rect 2196 21190 2206 21242
rect 2206 21190 2252 21242
rect 1956 21188 2012 21190
rect 2036 21188 2092 21190
rect 2116 21188 2172 21190
rect 2196 21188 2252 21190
rect 6956 21242 7012 21244
rect 7036 21242 7092 21244
rect 7116 21242 7172 21244
rect 7196 21242 7252 21244
rect 6956 21190 7002 21242
rect 7002 21190 7012 21242
rect 7036 21190 7066 21242
rect 7066 21190 7078 21242
rect 7078 21190 7092 21242
rect 7116 21190 7130 21242
rect 7130 21190 7142 21242
rect 7142 21190 7172 21242
rect 7196 21190 7206 21242
rect 7206 21190 7252 21242
rect 6956 21188 7012 21190
rect 7036 21188 7092 21190
rect 7116 21188 7172 21190
rect 7196 21188 7252 21190
rect 11956 21242 12012 21244
rect 12036 21242 12092 21244
rect 12116 21242 12172 21244
rect 12196 21242 12252 21244
rect 11956 21190 12002 21242
rect 12002 21190 12012 21242
rect 12036 21190 12066 21242
rect 12066 21190 12078 21242
rect 12078 21190 12092 21242
rect 12116 21190 12130 21242
rect 12130 21190 12142 21242
rect 12142 21190 12172 21242
rect 12196 21190 12206 21242
rect 12206 21190 12252 21242
rect 11956 21188 12012 21190
rect 12036 21188 12092 21190
rect 12116 21188 12172 21190
rect 12196 21188 12252 21190
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 17002 21242
rect 17002 21190 17012 21242
rect 17036 21190 17066 21242
rect 17066 21190 17078 21242
rect 17078 21190 17092 21242
rect 17116 21190 17130 21242
rect 17130 21190 17142 21242
rect 17142 21190 17172 21242
rect 17196 21190 17206 21242
rect 17206 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 2616 20698 2672 20700
rect 2696 20698 2752 20700
rect 2776 20698 2832 20700
rect 2856 20698 2912 20700
rect 2616 20646 2662 20698
rect 2662 20646 2672 20698
rect 2696 20646 2726 20698
rect 2726 20646 2738 20698
rect 2738 20646 2752 20698
rect 2776 20646 2790 20698
rect 2790 20646 2802 20698
rect 2802 20646 2832 20698
rect 2856 20646 2866 20698
rect 2866 20646 2912 20698
rect 2616 20644 2672 20646
rect 2696 20644 2752 20646
rect 2776 20644 2832 20646
rect 2856 20644 2912 20646
rect 7616 20698 7672 20700
rect 7696 20698 7752 20700
rect 7776 20698 7832 20700
rect 7856 20698 7912 20700
rect 7616 20646 7662 20698
rect 7662 20646 7672 20698
rect 7696 20646 7726 20698
rect 7726 20646 7738 20698
rect 7738 20646 7752 20698
rect 7776 20646 7790 20698
rect 7790 20646 7802 20698
rect 7802 20646 7832 20698
rect 7856 20646 7866 20698
rect 7866 20646 7912 20698
rect 7616 20644 7672 20646
rect 7696 20644 7752 20646
rect 7776 20644 7832 20646
rect 7856 20644 7912 20646
rect 12616 20698 12672 20700
rect 12696 20698 12752 20700
rect 12776 20698 12832 20700
rect 12856 20698 12912 20700
rect 12616 20646 12662 20698
rect 12662 20646 12672 20698
rect 12696 20646 12726 20698
rect 12726 20646 12738 20698
rect 12738 20646 12752 20698
rect 12776 20646 12790 20698
rect 12790 20646 12802 20698
rect 12802 20646 12832 20698
rect 12856 20646 12866 20698
rect 12866 20646 12912 20698
rect 12616 20644 12672 20646
rect 12696 20644 12752 20646
rect 12776 20644 12832 20646
rect 12856 20644 12912 20646
rect 1398 20576 1454 20632
rect 1956 20154 2012 20156
rect 2036 20154 2092 20156
rect 2116 20154 2172 20156
rect 2196 20154 2252 20156
rect 1956 20102 2002 20154
rect 2002 20102 2012 20154
rect 2036 20102 2066 20154
rect 2066 20102 2078 20154
rect 2078 20102 2092 20154
rect 2116 20102 2130 20154
rect 2130 20102 2142 20154
rect 2142 20102 2172 20154
rect 2196 20102 2206 20154
rect 2206 20102 2252 20154
rect 1956 20100 2012 20102
rect 2036 20100 2092 20102
rect 2116 20100 2172 20102
rect 2196 20100 2252 20102
rect 6956 20154 7012 20156
rect 7036 20154 7092 20156
rect 7116 20154 7172 20156
rect 7196 20154 7252 20156
rect 6956 20102 7002 20154
rect 7002 20102 7012 20154
rect 7036 20102 7066 20154
rect 7066 20102 7078 20154
rect 7078 20102 7092 20154
rect 7116 20102 7130 20154
rect 7130 20102 7142 20154
rect 7142 20102 7172 20154
rect 7196 20102 7206 20154
rect 7206 20102 7252 20154
rect 6956 20100 7012 20102
rect 7036 20100 7092 20102
rect 7116 20100 7172 20102
rect 7196 20100 7252 20102
rect 11956 20154 12012 20156
rect 12036 20154 12092 20156
rect 12116 20154 12172 20156
rect 12196 20154 12252 20156
rect 11956 20102 12002 20154
rect 12002 20102 12012 20154
rect 12036 20102 12066 20154
rect 12066 20102 12078 20154
rect 12078 20102 12092 20154
rect 12116 20102 12130 20154
rect 12130 20102 12142 20154
rect 12142 20102 12172 20154
rect 12196 20102 12206 20154
rect 12206 20102 12252 20154
rect 11956 20100 12012 20102
rect 12036 20100 12092 20102
rect 12116 20100 12172 20102
rect 12196 20100 12252 20102
rect 17616 20698 17672 20700
rect 17696 20698 17752 20700
rect 17776 20698 17832 20700
rect 17856 20698 17912 20700
rect 17616 20646 17662 20698
rect 17662 20646 17672 20698
rect 17696 20646 17726 20698
rect 17726 20646 17738 20698
rect 17738 20646 17752 20698
rect 17776 20646 17790 20698
rect 17790 20646 17802 20698
rect 17802 20646 17832 20698
rect 17856 20646 17866 20698
rect 17866 20646 17912 20698
rect 17616 20644 17672 20646
rect 17696 20644 17752 20646
rect 17776 20644 17832 20646
rect 17856 20644 17912 20646
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 17002 20154
rect 17002 20102 17012 20154
rect 17036 20102 17066 20154
rect 17066 20102 17078 20154
rect 17078 20102 17092 20154
rect 17116 20102 17130 20154
rect 17130 20102 17142 20154
rect 17142 20102 17172 20154
rect 17196 20102 17206 20154
rect 17206 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 938 19796 940 19816
rect 940 19796 992 19816
rect 992 19796 994 19816
rect 938 19760 994 19796
rect 2616 19610 2672 19612
rect 2696 19610 2752 19612
rect 2776 19610 2832 19612
rect 2856 19610 2912 19612
rect 2616 19558 2662 19610
rect 2662 19558 2672 19610
rect 2696 19558 2726 19610
rect 2726 19558 2738 19610
rect 2738 19558 2752 19610
rect 2776 19558 2790 19610
rect 2790 19558 2802 19610
rect 2802 19558 2832 19610
rect 2856 19558 2866 19610
rect 2866 19558 2912 19610
rect 2616 19556 2672 19558
rect 2696 19556 2752 19558
rect 2776 19556 2832 19558
rect 2856 19556 2912 19558
rect 7616 19610 7672 19612
rect 7696 19610 7752 19612
rect 7776 19610 7832 19612
rect 7856 19610 7912 19612
rect 7616 19558 7662 19610
rect 7662 19558 7672 19610
rect 7696 19558 7726 19610
rect 7726 19558 7738 19610
rect 7738 19558 7752 19610
rect 7776 19558 7790 19610
rect 7790 19558 7802 19610
rect 7802 19558 7832 19610
rect 7856 19558 7866 19610
rect 7866 19558 7912 19610
rect 7616 19556 7672 19558
rect 7696 19556 7752 19558
rect 7776 19556 7832 19558
rect 7856 19556 7912 19558
rect 12616 19610 12672 19612
rect 12696 19610 12752 19612
rect 12776 19610 12832 19612
rect 12856 19610 12912 19612
rect 12616 19558 12662 19610
rect 12662 19558 12672 19610
rect 12696 19558 12726 19610
rect 12726 19558 12738 19610
rect 12738 19558 12752 19610
rect 12776 19558 12790 19610
rect 12790 19558 12802 19610
rect 12802 19558 12832 19610
rect 12856 19558 12866 19610
rect 12866 19558 12912 19610
rect 12616 19556 12672 19558
rect 12696 19556 12752 19558
rect 12776 19556 12832 19558
rect 12856 19556 12912 19558
rect 17616 19610 17672 19612
rect 17696 19610 17752 19612
rect 17776 19610 17832 19612
rect 17856 19610 17912 19612
rect 17616 19558 17662 19610
rect 17662 19558 17672 19610
rect 17696 19558 17726 19610
rect 17726 19558 17738 19610
rect 17738 19558 17752 19610
rect 17776 19558 17790 19610
rect 17790 19558 17802 19610
rect 17802 19558 17832 19610
rect 17856 19558 17866 19610
rect 17866 19558 17912 19610
rect 17616 19556 17672 19558
rect 17696 19556 17752 19558
rect 17776 19556 17832 19558
rect 17856 19556 17912 19558
rect 1398 19116 1400 19136
rect 1400 19116 1452 19136
rect 1452 19116 1454 19136
rect 1398 19080 1454 19116
rect 1956 19066 2012 19068
rect 2036 19066 2092 19068
rect 2116 19066 2172 19068
rect 2196 19066 2252 19068
rect 1956 19014 2002 19066
rect 2002 19014 2012 19066
rect 2036 19014 2066 19066
rect 2066 19014 2078 19066
rect 2078 19014 2092 19066
rect 2116 19014 2130 19066
rect 2130 19014 2142 19066
rect 2142 19014 2172 19066
rect 2196 19014 2206 19066
rect 2206 19014 2252 19066
rect 1956 19012 2012 19014
rect 2036 19012 2092 19014
rect 2116 19012 2172 19014
rect 2196 19012 2252 19014
rect 6956 19066 7012 19068
rect 7036 19066 7092 19068
rect 7116 19066 7172 19068
rect 7196 19066 7252 19068
rect 6956 19014 7002 19066
rect 7002 19014 7012 19066
rect 7036 19014 7066 19066
rect 7066 19014 7078 19066
rect 7078 19014 7092 19066
rect 7116 19014 7130 19066
rect 7130 19014 7142 19066
rect 7142 19014 7172 19066
rect 7196 19014 7206 19066
rect 7206 19014 7252 19066
rect 6956 19012 7012 19014
rect 7036 19012 7092 19014
rect 7116 19012 7172 19014
rect 7196 19012 7252 19014
rect 11956 19066 12012 19068
rect 12036 19066 12092 19068
rect 12116 19066 12172 19068
rect 12196 19066 12252 19068
rect 11956 19014 12002 19066
rect 12002 19014 12012 19066
rect 12036 19014 12066 19066
rect 12066 19014 12078 19066
rect 12078 19014 12092 19066
rect 12116 19014 12130 19066
rect 12130 19014 12142 19066
rect 12142 19014 12172 19066
rect 12196 19014 12206 19066
rect 12206 19014 12252 19066
rect 11956 19012 12012 19014
rect 12036 19012 12092 19014
rect 12116 19012 12172 19014
rect 12196 19012 12252 19014
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 17002 19066
rect 17002 19014 17012 19066
rect 17036 19014 17066 19066
rect 17066 19014 17078 19066
rect 17078 19014 17092 19066
rect 17116 19014 17130 19066
rect 17130 19014 17142 19066
rect 17142 19014 17172 19066
rect 17196 19014 17206 19066
rect 17206 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 18970 19352 19026 19408
rect 2616 18522 2672 18524
rect 2696 18522 2752 18524
rect 2776 18522 2832 18524
rect 2856 18522 2912 18524
rect 2616 18470 2662 18522
rect 2662 18470 2672 18522
rect 2696 18470 2726 18522
rect 2726 18470 2738 18522
rect 2738 18470 2752 18522
rect 2776 18470 2790 18522
rect 2790 18470 2802 18522
rect 2802 18470 2832 18522
rect 2856 18470 2866 18522
rect 2866 18470 2912 18522
rect 2616 18468 2672 18470
rect 2696 18468 2752 18470
rect 2776 18468 2832 18470
rect 2856 18468 2912 18470
rect 7616 18522 7672 18524
rect 7696 18522 7752 18524
rect 7776 18522 7832 18524
rect 7856 18522 7912 18524
rect 7616 18470 7662 18522
rect 7662 18470 7672 18522
rect 7696 18470 7726 18522
rect 7726 18470 7738 18522
rect 7738 18470 7752 18522
rect 7776 18470 7790 18522
rect 7790 18470 7802 18522
rect 7802 18470 7832 18522
rect 7856 18470 7866 18522
rect 7866 18470 7912 18522
rect 7616 18468 7672 18470
rect 7696 18468 7752 18470
rect 7776 18468 7832 18470
rect 7856 18468 7912 18470
rect 12616 18522 12672 18524
rect 12696 18522 12752 18524
rect 12776 18522 12832 18524
rect 12856 18522 12912 18524
rect 12616 18470 12662 18522
rect 12662 18470 12672 18522
rect 12696 18470 12726 18522
rect 12726 18470 12738 18522
rect 12738 18470 12752 18522
rect 12776 18470 12790 18522
rect 12790 18470 12802 18522
rect 12802 18470 12832 18522
rect 12856 18470 12866 18522
rect 12866 18470 12912 18522
rect 12616 18468 12672 18470
rect 12696 18468 12752 18470
rect 12776 18468 12832 18470
rect 12856 18468 12912 18470
rect 17616 18522 17672 18524
rect 17696 18522 17752 18524
rect 17776 18522 17832 18524
rect 17856 18522 17912 18524
rect 17616 18470 17662 18522
rect 17662 18470 17672 18522
rect 17696 18470 17726 18522
rect 17726 18470 17738 18522
rect 17738 18470 17752 18522
rect 17776 18470 17790 18522
rect 17790 18470 17802 18522
rect 17802 18470 17832 18522
rect 17856 18470 17866 18522
rect 17866 18470 17912 18522
rect 17616 18468 17672 18470
rect 17696 18468 17752 18470
rect 17776 18468 17832 18470
rect 17856 18468 17912 18470
rect 938 18400 994 18456
rect 21956 21242 22012 21244
rect 22036 21242 22092 21244
rect 22116 21242 22172 21244
rect 22196 21242 22252 21244
rect 21956 21190 22002 21242
rect 22002 21190 22012 21242
rect 22036 21190 22066 21242
rect 22066 21190 22078 21242
rect 22078 21190 22092 21242
rect 22116 21190 22130 21242
rect 22130 21190 22142 21242
rect 22142 21190 22172 21242
rect 22196 21190 22206 21242
rect 22206 21190 22252 21242
rect 21956 21188 22012 21190
rect 22036 21188 22092 21190
rect 22116 21188 22172 21190
rect 22196 21188 22252 21190
rect 26956 21242 27012 21244
rect 27036 21242 27092 21244
rect 27116 21242 27172 21244
rect 27196 21242 27252 21244
rect 26956 21190 27002 21242
rect 27002 21190 27012 21242
rect 27036 21190 27066 21242
rect 27066 21190 27078 21242
rect 27078 21190 27092 21242
rect 27116 21190 27130 21242
rect 27130 21190 27142 21242
rect 27142 21190 27172 21242
rect 27196 21190 27206 21242
rect 27206 21190 27252 21242
rect 26956 21188 27012 21190
rect 27036 21188 27092 21190
rect 27116 21188 27172 21190
rect 27196 21188 27252 21190
rect 31956 21242 32012 21244
rect 32036 21242 32092 21244
rect 32116 21242 32172 21244
rect 32196 21242 32252 21244
rect 31956 21190 32002 21242
rect 32002 21190 32012 21242
rect 32036 21190 32066 21242
rect 32066 21190 32078 21242
rect 32078 21190 32092 21242
rect 32116 21190 32130 21242
rect 32130 21190 32142 21242
rect 32142 21190 32172 21242
rect 32196 21190 32206 21242
rect 32206 21190 32252 21242
rect 31956 21188 32012 21190
rect 32036 21188 32092 21190
rect 32116 21188 32172 21190
rect 32196 21188 32252 21190
rect 36956 21242 37012 21244
rect 37036 21242 37092 21244
rect 37116 21242 37172 21244
rect 37196 21242 37252 21244
rect 36956 21190 37002 21242
rect 37002 21190 37012 21242
rect 37036 21190 37066 21242
rect 37066 21190 37078 21242
rect 37078 21190 37092 21242
rect 37116 21190 37130 21242
rect 37130 21190 37142 21242
rect 37142 21190 37172 21242
rect 37196 21190 37206 21242
rect 37206 21190 37252 21242
rect 36956 21188 37012 21190
rect 37036 21188 37092 21190
rect 37116 21188 37172 21190
rect 37196 21188 37252 21190
rect 22616 20698 22672 20700
rect 22696 20698 22752 20700
rect 22776 20698 22832 20700
rect 22856 20698 22912 20700
rect 22616 20646 22662 20698
rect 22662 20646 22672 20698
rect 22696 20646 22726 20698
rect 22726 20646 22738 20698
rect 22738 20646 22752 20698
rect 22776 20646 22790 20698
rect 22790 20646 22802 20698
rect 22802 20646 22832 20698
rect 22856 20646 22866 20698
rect 22866 20646 22912 20698
rect 22616 20644 22672 20646
rect 22696 20644 22752 20646
rect 22776 20644 22832 20646
rect 22856 20644 22912 20646
rect 27616 20698 27672 20700
rect 27696 20698 27752 20700
rect 27776 20698 27832 20700
rect 27856 20698 27912 20700
rect 27616 20646 27662 20698
rect 27662 20646 27672 20698
rect 27696 20646 27726 20698
rect 27726 20646 27738 20698
rect 27738 20646 27752 20698
rect 27776 20646 27790 20698
rect 27790 20646 27802 20698
rect 27802 20646 27832 20698
rect 27856 20646 27866 20698
rect 27866 20646 27912 20698
rect 27616 20644 27672 20646
rect 27696 20644 27752 20646
rect 27776 20644 27832 20646
rect 27856 20644 27912 20646
rect 32616 20698 32672 20700
rect 32696 20698 32752 20700
rect 32776 20698 32832 20700
rect 32856 20698 32912 20700
rect 32616 20646 32662 20698
rect 32662 20646 32672 20698
rect 32696 20646 32726 20698
rect 32726 20646 32738 20698
rect 32738 20646 32752 20698
rect 32776 20646 32790 20698
rect 32790 20646 32802 20698
rect 32802 20646 32832 20698
rect 32856 20646 32866 20698
rect 32866 20646 32912 20698
rect 32616 20644 32672 20646
rect 32696 20644 32752 20646
rect 32776 20644 32832 20646
rect 32856 20644 32912 20646
rect 21956 20154 22012 20156
rect 22036 20154 22092 20156
rect 22116 20154 22172 20156
rect 22196 20154 22252 20156
rect 21956 20102 22002 20154
rect 22002 20102 22012 20154
rect 22036 20102 22066 20154
rect 22066 20102 22078 20154
rect 22078 20102 22092 20154
rect 22116 20102 22130 20154
rect 22130 20102 22142 20154
rect 22142 20102 22172 20154
rect 22196 20102 22206 20154
rect 22206 20102 22252 20154
rect 21956 20100 22012 20102
rect 22036 20100 22092 20102
rect 22116 20100 22172 20102
rect 22196 20100 22252 20102
rect 26956 20154 27012 20156
rect 27036 20154 27092 20156
rect 27116 20154 27172 20156
rect 27196 20154 27252 20156
rect 26956 20102 27002 20154
rect 27002 20102 27012 20154
rect 27036 20102 27066 20154
rect 27066 20102 27078 20154
rect 27078 20102 27092 20154
rect 27116 20102 27130 20154
rect 27130 20102 27142 20154
rect 27142 20102 27172 20154
rect 27196 20102 27206 20154
rect 27206 20102 27252 20154
rect 26956 20100 27012 20102
rect 27036 20100 27092 20102
rect 27116 20100 27172 20102
rect 27196 20100 27252 20102
rect 31956 20154 32012 20156
rect 32036 20154 32092 20156
rect 32116 20154 32172 20156
rect 32196 20154 32252 20156
rect 31956 20102 32002 20154
rect 32002 20102 32012 20154
rect 32036 20102 32066 20154
rect 32066 20102 32078 20154
rect 32078 20102 32092 20154
rect 32116 20102 32130 20154
rect 32130 20102 32142 20154
rect 32142 20102 32172 20154
rect 32196 20102 32206 20154
rect 32206 20102 32252 20154
rect 31956 20100 32012 20102
rect 32036 20100 32092 20102
rect 32116 20100 32172 20102
rect 32196 20100 32252 20102
rect 38474 21836 38476 21856
rect 38476 21836 38528 21856
rect 38528 21836 38530 21856
rect 38474 21800 38530 21836
rect 37616 21786 37672 21788
rect 37696 21786 37752 21788
rect 37776 21786 37832 21788
rect 37856 21786 37912 21788
rect 37616 21734 37662 21786
rect 37662 21734 37672 21786
rect 37696 21734 37726 21786
rect 37726 21734 37738 21786
rect 37738 21734 37752 21786
rect 37776 21734 37790 21786
rect 37790 21734 37802 21786
rect 37802 21734 37832 21786
rect 37856 21734 37866 21786
rect 37866 21734 37912 21786
rect 37616 21732 37672 21734
rect 37696 21732 37752 21734
rect 37776 21732 37832 21734
rect 37856 21732 37912 21734
rect 37616 20698 37672 20700
rect 37696 20698 37752 20700
rect 37776 20698 37832 20700
rect 37856 20698 37912 20700
rect 37616 20646 37662 20698
rect 37662 20646 37672 20698
rect 37696 20646 37726 20698
rect 37726 20646 37738 20698
rect 37738 20646 37752 20698
rect 37776 20646 37790 20698
rect 37790 20646 37802 20698
rect 37802 20646 37832 20698
rect 37856 20646 37866 20698
rect 37866 20646 37912 20698
rect 37616 20644 37672 20646
rect 37696 20644 37752 20646
rect 37776 20644 37832 20646
rect 37856 20644 37912 20646
rect 38474 21120 38530 21176
rect 39026 20440 39082 20496
rect 36956 20154 37012 20156
rect 37036 20154 37092 20156
rect 37116 20154 37172 20156
rect 37196 20154 37252 20156
rect 36956 20102 37002 20154
rect 37002 20102 37012 20154
rect 37036 20102 37066 20154
rect 37066 20102 37078 20154
rect 37078 20102 37092 20154
rect 37116 20102 37130 20154
rect 37130 20102 37142 20154
rect 37142 20102 37172 20154
rect 37196 20102 37206 20154
rect 37206 20102 37252 20154
rect 36956 20100 37012 20102
rect 37036 20100 37092 20102
rect 37116 20100 37172 20102
rect 37196 20100 37252 20102
rect 21956 19066 22012 19068
rect 22036 19066 22092 19068
rect 22116 19066 22172 19068
rect 22196 19066 22252 19068
rect 21956 19014 22002 19066
rect 22002 19014 22012 19066
rect 22036 19014 22066 19066
rect 22066 19014 22078 19066
rect 22078 19014 22092 19066
rect 22116 19014 22130 19066
rect 22130 19014 22142 19066
rect 22142 19014 22172 19066
rect 22196 19014 22206 19066
rect 22206 19014 22252 19066
rect 21956 19012 22012 19014
rect 22036 19012 22092 19014
rect 22116 19012 22172 19014
rect 22196 19012 22252 19014
rect 22616 19610 22672 19612
rect 22696 19610 22752 19612
rect 22776 19610 22832 19612
rect 22856 19610 22912 19612
rect 22616 19558 22662 19610
rect 22662 19558 22672 19610
rect 22696 19558 22726 19610
rect 22726 19558 22738 19610
rect 22738 19558 22752 19610
rect 22776 19558 22790 19610
rect 22790 19558 22802 19610
rect 22802 19558 22832 19610
rect 22856 19558 22866 19610
rect 22866 19558 22912 19610
rect 22616 19556 22672 19558
rect 22696 19556 22752 19558
rect 22776 19556 22832 19558
rect 22856 19556 22912 19558
rect 38842 19760 38898 19816
rect 27616 19610 27672 19612
rect 27696 19610 27752 19612
rect 27776 19610 27832 19612
rect 27856 19610 27912 19612
rect 27616 19558 27662 19610
rect 27662 19558 27672 19610
rect 27696 19558 27726 19610
rect 27726 19558 27738 19610
rect 27738 19558 27752 19610
rect 27776 19558 27790 19610
rect 27790 19558 27802 19610
rect 27802 19558 27832 19610
rect 27856 19558 27866 19610
rect 27866 19558 27912 19610
rect 27616 19556 27672 19558
rect 27696 19556 27752 19558
rect 27776 19556 27832 19558
rect 27856 19556 27912 19558
rect 32616 19610 32672 19612
rect 32696 19610 32752 19612
rect 32776 19610 32832 19612
rect 32856 19610 32912 19612
rect 32616 19558 32662 19610
rect 32662 19558 32672 19610
rect 32696 19558 32726 19610
rect 32726 19558 32738 19610
rect 32738 19558 32752 19610
rect 32776 19558 32790 19610
rect 32790 19558 32802 19610
rect 32802 19558 32832 19610
rect 32856 19558 32866 19610
rect 32866 19558 32912 19610
rect 32616 19556 32672 19558
rect 32696 19556 32752 19558
rect 32776 19556 32832 19558
rect 32856 19556 32912 19558
rect 26956 19066 27012 19068
rect 27036 19066 27092 19068
rect 27116 19066 27172 19068
rect 27196 19066 27252 19068
rect 26956 19014 27002 19066
rect 27002 19014 27012 19066
rect 27036 19014 27066 19066
rect 27066 19014 27078 19066
rect 27078 19014 27092 19066
rect 27116 19014 27130 19066
rect 27130 19014 27142 19066
rect 27142 19014 27172 19066
rect 27196 19014 27206 19066
rect 27206 19014 27252 19066
rect 26956 19012 27012 19014
rect 27036 19012 27092 19014
rect 27116 19012 27172 19014
rect 27196 19012 27252 19014
rect 22616 18522 22672 18524
rect 22696 18522 22752 18524
rect 22776 18522 22832 18524
rect 22856 18522 22912 18524
rect 22616 18470 22662 18522
rect 22662 18470 22672 18522
rect 22696 18470 22726 18522
rect 22726 18470 22738 18522
rect 22738 18470 22752 18522
rect 22776 18470 22790 18522
rect 22790 18470 22802 18522
rect 22802 18470 22832 18522
rect 22856 18470 22866 18522
rect 22866 18470 22912 18522
rect 22616 18468 22672 18470
rect 22696 18468 22752 18470
rect 22776 18468 22832 18470
rect 22856 18468 22912 18470
rect 27616 18522 27672 18524
rect 27696 18522 27752 18524
rect 27776 18522 27832 18524
rect 27856 18522 27912 18524
rect 27616 18470 27662 18522
rect 27662 18470 27672 18522
rect 27696 18470 27726 18522
rect 27726 18470 27738 18522
rect 27738 18470 27752 18522
rect 27776 18470 27790 18522
rect 27790 18470 27802 18522
rect 27802 18470 27832 18522
rect 27856 18470 27866 18522
rect 27866 18470 27912 18522
rect 27616 18468 27672 18470
rect 27696 18468 27752 18470
rect 27776 18468 27832 18470
rect 27856 18468 27912 18470
rect 1956 17978 2012 17980
rect 2036 17978 2092 17980
rect 2116 17978 2172 17980
rect 2196 17978 2252 17980
rect 1956 17926 2002 17978
rect 2002 17926 2012 17978
rect 2036 17926 2066 17978
rect 2066 17926 2078 17978
rect 2078 17926 2092 17978
rect 2116 17926 2130 17978
rect 2130 17926 2142 17978
rect 2142 17926 2172 17978
rect 2196 17926 2206 17978
rect 2206 17926 2252 17978
rect 1956 17924 2012 17926
rect 2036 17924 2092 17926
rect 2116 17924 2172 17926
rect 2196 17924 2252 17926
rect 6956 17978 7012 17980
rect 7036 17978 7092 17980
rect 7116 17978 7172 17980
rect 7196 17978 7252 17980
rect 6956 17926 7002 17978
rect 7002 17926 7012 17978
rect 7036 17926 7066 17978
rect 7066 17926 7078 17978
rect 7078 17926 7092 17978
rect 7116 17926 7130 17978
rect 7130 17926 7142 17978
rect 7142 17926 7172 17978
rect 7196 17926 7206 17978
rect 7206 17926 7252 17978
rect 6956 17924 7012 17926
rect 7036 17924 7092 17926
rect 7116 17924 7172 17926
rect 7196 17924 7252 17926
rect 11956 17978 12012 17980
rect 12036 17978 12092 17980
rect 12116 17978 12172 17980
rect 12196 17978 12252 17980
rect 11956 17926 12002 17978
rect 12002 17926 12012 17978
rect 12036 17926 12066 17978
rect 12066 17926 12078 17978
rect 12078 17926 12092 17978
rect 12116 17926 12130 17978
rect 12130 17926 12142 17978
rect 12142 17926 12172 17978
rect 12196 17926 12206 17978
rect 12206 17926 12252 17978
rect 11956 17924 12012 17926
rect 12036 17924 12092 17926
rect 12116 17924 12172 17926
rect 12196 17924 12252 17926
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 17002 17978
rect 17002 17926 17012 17978
rect 17036 17926 17066 17978
rect 17066 17926 17078 17978
rect 17078 17926 17092 17978
rect 17116 17926 17130 17978
rect 17130 17926 17142 17978
rect 17142 17926 17172 17978
rect 17196 17926 17206 17978
rect 17206 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 21956 17978 22012 17980
rect 22036 17978 22092 17980
rect 22116 17978 22172 17980
rect 22196 17978 22252 17980
rect 21956 17926 22002 17978
rect 22002 17926 22012 17978
rect 22036 17926 22066 17978
rect 22066 17926 22078 17978
rect 22078 17926 22092 17978
rect 22116 17926 22130 17978
rect 22130 17926 22142 17978
rect 22142 17926 22172 17978
rect 22196 17926 22206 17978
rect 22206 17926 22252 17978
rect 21956 17924 22012 17926
rect 22036 17924 22092 17926
rect 22116 17924 22172 17926
rect 22196 17924 22252 17926
rect 26956 17978 27012 17980
rect 27036 17978 27092 17980
rect 27116 17978 27172 17980
rect 27196 17978 27252 17980
rect 26956 17926 27002 17978
rect 27002 17926 27012 17978
rect 27036 17926 27066 17978
rect 27066 17926 27078 17978
rect 27078 17926 27092 17978
rect 27116 17926 27130 17978
rect 27130 17926 27142 17978
rect 27142 17926 27172 17978
rect 27196 17926 27206 17978
rect 27206 17926 27252 17978
rect 26956 17924 27012 17926
rect 27036 17924 27092 17926
rect 27116 17924 27172 17926
rect 27196 17924 27252 17926
rect 31956 19066 32012 19068
rect 32036 19066 32092 19068
rect 32116 19066 32172 19068
rect 32196 19066 32252 19068
rect 31956 19014 32002 19066
rect 32002 19014 32012 19066
rect 32036 19014 32066 19066
rect 32066 19014 32078 19066
rect 32078 19014 32092 19066
rect 32116 19014 32130 19066
rect 32130 19014 32142 19066
rect 32142 19014 32172 19066
rect 32196 19014 32206 19066
rect 32206 19014 32252 19066
rect 31956 19012 32012 19014
rect 32036 19012 32092 19014
rect 32116 19012 32172 19014
rect 32196 19012 32252 19014
rect 36956 19066 37012 19068
rect 37036 19066 37092 19068
rect 37116 19066 37172 19068
rect 37196 19066 37252 19068
rect 36956 19014 37002 19066
rect 37002 19014 37012 19066
rect 37036 19014 37066 19066
rect 37066 19014 37078 19066
rect 37078 19014 37092 19066
rect 37116 19014 37130 19066
rect 37130 19014 37142 19066
rect 37142 19014 37172 19066
rect 37196 19014 37206 19066
rect 37206 19014 37252 19066
rect 36956 19012 37012 19014
rect 37036 19012 37092 19014
rect 37116 19012 37172 19014
rect 37196 19012 37252 19014
rect 37616 19610 37672 19612
rect 37696 19610 37752 19612
rect 37776 19610 37832 19612
rect 37856 19610 37912 19612
rect 37616 19558 37662 19610
rect 37662 19558 37672 19610
rect 37696 19558 37726 19610
rect 37726 19558 37738 19610
rect 37738 19558 37752 19610
rect 37776 19558 37790 19610
rect 37790 19558 37802 19610
rect 37802 19558 37832 19610
rect 37856 19558 37866 19610
rect 37866 19558 37912 19610
rect 37616 19556 37672 19558
rect 37696 19556 37752 19558
rect 37776 19556 37832 19558
rect 37856 19556 37912 19558
rect 38290 19372 38346 19408
rect 38290 19352 38292 19372
rect 38292 19352 38344 19372
rect 38344 19352 38346 19372
rect 38474 19116 38476 19136
rect 38476 19116 38528 19136
rect 38528 19116 38530 19136
rect 38474 19080 38530 19116
rect 32616 18522 32672 18524
rect 32696 18522 32752 18524
rect 32776 18522 32832 18524
rect 32856 18522 32912 18524
rect 32616 18470 32662 18522
rect 32662 18470 32672 18522
rect 32696 18470 32726 18522
rect 32726 18470 32738 18522
rect 32738 18470 32752 18522
rect 32776 18470 32790 18522
rect 32790 18470 32802 18522
rect 32802 18470 32832 18522
rect 32856 18470 32866 18522
rect 32866 18470 32912 18522
rect 32616 18468 32672 18470
rect 32696 18468 32752 18470
rect 32776 18468 32832 18470
rect 32856 18468 32912 18470
rect 37616 18522 37672 18524
rect 37696 18522 37752 18524
rect 37776 18522 37832 18524
rect 37856 18522 37912 18524
rect 37616 18470 37662 18522
rect 37662 18470 37672 18522
rect 37696 18470 37726 18522
rect 37726 18470 37738 18522
rect 37738 18470 37752 18522
rect 37776 18470 37790 18522
rect 37790 18470 37802 18522
rect 37802 18470 37832 18522
rect 37856 18470 37866 18522
rect 37866 18470 37912 18522
rect 37616 18468 37672 18470
rect 37696 18468 37752 18470
rect 37776 18468 37832 18470
rect 37856 18468 37912 18470
rect 38474 18400 38530 18456
rect 31956 17978 32012 17980
rect 32036 17978 32092 17980
rect 32116 17978 32172 17980
rect 32196 17978 32252 17980
rect 31956 17926 32002 17978
rect 32002 17926 32012 17978
rect 32036 17926 32066 17978
rect 32066 17926 32078 17978
rect 32078 17926 32092 17978
rect 32116 17926 32130 17978
rect 32130 17926 32142 17978
rect 32142 17926 32172 17978
rect 32196 17926 32206 17978
rect 32206 17926 32252 17978
rect 31956 17924 32012 17926
rect 32036 17924 32092 17926
rect 32116 17924 32172 17926
rect 32196 17924 32252 17926
rect 36956 17978 37012 17980
rect 37036 17978 37092 17980
rect 37116 17978 37172 17980
rect 37196 17978 37252 17980
rect 36956 17926 37002 17978
rect 37002 17926 37012 17978
rect 37036 17926 37066 17978
rect 37066 17926 37078 17978
rect 37078 17926 37092 17978
rect 37116 17926 37130 17978
rect 37130 17926 37142 17978
rect 37142 17926 37172 17978
rect 37196 17926 37206 17978
rect 37206 17926 37252 17978
rect 36956 17924 37012 17926
rect 37036 17924 37092 17926
rect 37116 17924 37172 17926
rect 37196 17924 37252 17926
rect 34518 17720 34574 17776
rect 2616 17434 2672 17436
rect 2696 17434 2752 17436
rect 2776 17434 2832 17436
rect 2856 17434 2912 17436
rect 2616 17382 2662 17434
rect 2662 17382 2672 17434
rect 2696 17382 2726 17434
rect 2726 17382 2738 17434
rect 2738 17382 2752 17434
rect 2776 17382 2790 17434
rect 2790 17382 2802 17434
rect 2802 17382 2832 17434
rect 2856 17382 2866 17434
rect 2866 17382 2912 17434
rect 2616 17380 2672 17382
rect 2696 17380 2752 17382
rect 2776 17380 2832 17382
rect 2856 17380 2912 17382
rect 7616 17434 7672 17436
rect 7696 17434 7752 17436
rect 7776 17434 7832 17436
rect 7856 17434 7912 17436
rect 7616 17382 7662 17434
rect 7662 17382 7672 17434
rect 7696 17382 7726 17434
rect 7726 17382 7738 17434
rect 7738 17382 7752 17434
rect 7776 17382 7790 17434
rect 7790 17382 7802 17434
rect 7802 17382 7832 17434
rect 7856 17382 7866 17434
rect 7866 17382 7912 17434
rect 7616 17380 7672 17382
rect 7696 17380 7752 17382
rect 7776 17380 7832 17382
rect 7856 17380 7912 17382
rect 12616 17434 12672 17436
rect 12696 17434 12752 17436
rect 12776 17434 12832 17436
rect 12856 17434 12912 17436
rect 12616 17382 12662 17434
rect 12662 17382 12672 17434
rect 12696 17382 12726 17434
rect 12726 17382 12738 17434
rect 12738 17382 12752 17434
rect 12776 17382 12790 17434
rect 12790 17382 12802 17434
rect 12802 17382 12832 17434
rect 12856 17382 12866 17434
rect 12866 17382 12912 17434
rect 12616 17380 12672 17382
rect 12696 17380 12752 17382
rect 12776 17380 12832 17382
rect 12856 17380 12912 17382
rect 17616 17434 17672 17436
rect 17696 17434 17752 17436
rect 17776 17434 17832 17436
rect 17856 17434 17912 17436
rect 17616 17382 17662 17434
rect 17662 17382 17672 17434
rect 17696 17382 17726 17434
rect 17726 17382 17738 17434
rect 17738 17382 17752 17434
rect 17776 17382 17790 17434
rect 17790 17382 17802 17434
rect 17802 17382 17832 17434
rect 17856 17382 17866 17434
rect 17866 17382 17912 17434
rect 17616 17380 17672 17382
rect 17696 17380 17752 17382
rect 17776 17380 17832 17382
rect 17856 17380 17912 17382
rect 22616 17434 22672 17436
rect 22696 17434 22752 17436
rect 22776 17434 22832 17436
rect 22856 17434 22912 17436
rect 22616 17382 22662 17434
rect 22662 17382 22672 17434
rect 22696 17382 22726 17434
rect 22726 17382 22738 17434
rect 22738 17382 22752 17434
rect 22776 17382 22790 17434
rect 22790 17382 22802 17434
rect 22802 17382 22832 17434
rect 22856 17382 22866 17434
rect 22866 17382 22912 17434
rect 22616 17380 22672 17382
rect 22696 17380 22752 17382
rect 22776 17380 22832 17382
rect 22856 17380 22912 17382
rect 27616 17434 27672 17436
rect 27696 17434 27752 17436
rect 27776 17434 27832 17436
rect 27856 17434 27912 17436
rect 27616 17382 27662 17434
rect 27662 17382 27672 17434
rect 27696 17382 27726 17434
rect 27726 17382 27738 17434
rect 27738 17382 27752 17434
rect 27776 17382 27790 17434
rect 27790 17382 27802 17434
rect 27802 17382 27832 17434
rect 27856 17382 27866 17434
rect 27866 17382 27912 17434
rect 27616 17380 27672 17382
rect 27696 17380 27752 17382
rect 27776 17380 27832 17382
rect 27856 17380 27912 17382
rect 32616 17434 32672 17436
rect 32696 17434 32752 17436
rect 32776 17434 32832 17436
rect 32856 17434 32912 17436
rect 32616 17382 32662 17434
rect 32662 17382 32672 17434
rect 32696 17382 32726 17434
rect 32726 17382 32738 17434
rect 32738 17382 32752 17434
rect 32776 17382 32790 17434
rect 32790 17382 32802 17434
rect 32802 17382 32832 17434
rect 32856 17382 32866 17434
rect 32866 17382 32912 17434
rect 32616 17380 32672 17382
rect 32696 17380 32752 17382
rect 32776 17380 32832 17382
rect 32856 17380 32912 17382
rect 37616 17434 37672 17436
rect 37696 17434 37752 17436
rect 37776 17434 37832 17436
rect 37856 17434 37912 17436
rect 37616 17382 37662 17434
rect 37662 17382 37672 17434
rect 37696 17382 37726 17434
rect 37726 17382 37738 17434
rect 37738 17382 37752 17434
rect 37776 17382 37790 17434
rect 37790 17382 37802 17434
rect 37802 17382 37832 17434
rect 37856 17382 37866 17434
rect 37866 17382 37912 17434
rect 37616 17380 37672 17382
rect 37696 17380 37752 17382
rect 37776 17380 37832 17382
rect 37856 17380 37912 17382
rect 1956 16890 2012 16892
rect 2036 16890 2092 16892
rect 2116 16890 2172 16892
rect 2196 16890 2252 16892
rect 1956 16838 2002 16890
rect 2002 16838 2012 16890
rect 2036 16838 2066 16890
rect 2066 16838 2078 16890
rect 2078 16838 2092 16890
rect 2116 16838 2130 16890
rect 2130 16838 2142 16890
rect 2142 16838 2172 16890
rect 2196 16838 2206 16890
rect 2206 16838 2252 16890
rect 1956 16836 2012 16838
rect 2036 16836 2092 16838
rect 2116 16836 2172 16838
rect 2196 16836 2252 16838
rect 6956 16890 7012 16892
rect 7036 16890 7092 16892
rect 7116 16890 7172 16892
rect 7196 16890 7252 16892
rect 6956 16838 7002 16890
rect 7002 16838 7012 16890
rect 7036 16838 7066 16890
rect 7066 16838 7078 16890
rect 7078 16838 7092 16890
rect 7116 16838 7130 16890
rect 7130 16838 7142 16890
rect 7142 16838 7172 16890
rect 7196 16838 7206 16890
rect 7206 16838 7252 16890
rect 6956 16836 7012 16838
rect 7036 16836 7092 16838
rect 7116 16836 7172 16838
rect 7196 16836 7252 16838
rect 11956 16890 12012 16892
rect 12036 16890 12092 16892
rect 12116 16890 12172 16892
rect 12196 16890 12252 16892
rect 11956 16838 12002 16890
rect 12002 16838 12012 16890
rect 12036 16838 12066 16890
rect 12066 16838 12078 16890
rect 12078 16838 12092 16890
rect 12116 16838 12130 16890
rect 12130 16838 12142 16890
rect 12142 16838 12172 16890
rect 12196 16838 12206 16890
rect 12206 16838 12252 16890
rect 11956 16836 12012 16838
rect 12036 16836 12092 16838
rect 12116 16836 12172 16838
rect 12196 16836 12252 16838
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 17002 16890
rect 17002 16838 17012 16890
rect 17036 16838 17066 16890
rect 17066 16838 17078 16890
rect 17078 16838 17092 16890
rect 17116 16838 17130 16890
rect 17130 16838 17142 16890
rect 17142 16838 17172 16890
rect 17196 16838 17206 16890
rect 17206 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 21956 16890 22012 16892
rect 22036 16890 22092 16892
rect 22116 16890 22172 16892
rect 22196 16890 22252 16892
rect 21956 16838 22002 16890
rect 22002 16838 22012 16890
rect 22036 16838 22066 16890
rect 22066 16838 22078 16890
rect 22078 16838 22092 16890
rect 22116 16838 22130 16890
rect 22130 16838 22142 16890
rect 22142 16838 22172 16890
rect 22196 16838 22206 16890
rect 22206 16838 22252 16890
rect 21956 16836 22012 16838
rect 22036 16836 22092 16838
rect 22116 16836 22172 16838
rect 22196 16836 22252 16838
rect 26956 16890 27012 16892
rect 27036 16890 27092 16892
rect 27116 16890 27172 16892
rect 27196 16890 27252 16892
rect 26956 16838 27002 16890
rect 27002 16838 27012 16890
rect 27036 16838 27066 16890
rect 27066 16838 27078 16890
rect 27078 16838 27092 16890
rect 27116 16838 27130 16890
rect 27130 16838 27142 16890
rect 27142 16838 27172 16890
rect 27196 16838 27206 16890
rect 27206 16838 27252 16890
rect 26956 16836 27012 16838
rect 27036 16836 27092 16838
rect 27116 16836 27172 16838
rect 27196 16836 27252 16838
rect 31956 16890 32012 16892
rect 32036 16890 32092 16892
rect 32116 16890 32172 16892
rect 32196 16890 32252 16892
rect 31956 16838 32002 16890
rect 32002 16838 32012 16890
rect 32036 16838 32066 16890
rect 32066 16838 32078 16890
rect 32078 16838 32092 16890
rect 32116 16838 32130 16890
rect 32130 16838 32142 16890
rect 32142 16838 32172 16890
rect 32196 16838 32206 16890
rect 32206 16838 32252 16890
rect 31956 16836 32012 16838
rect 32036 16836 32092 16838
rect 32116 16836 32172 16838
rect 32196 16836 32252 16838
rect 36956 16890 37012 16892
rect 37036 16890 37092 16892
rect 37116 16890 37172 16892
rect 37196 16890 37252 16892
rect 36956 16838 37002 16890
rect 37002 16838 37012 16890
rect 37036 16838 37066 16890
rect 37066 16838 37078 16890
rect 37078 16838 37092 16890
rect 37116 16838 37130 16890
rect 37130 16838 37142 16890
rect 37142 16838 37172 16890
rect 37196 16838 37206 16890
rect 37206 16838 37252 16890
rect 36956 16836 37012 16838
rect 37036 16836 37092 16838
rect 37116 16836 37172 16838
rect 37196 16836 37252 16838
rect 2616 16346 2672 16348
rect 2696 16346 2752 16348
rect 2776 16346 2832 16348
rect 2856 16346 2912 16348
rect 2616 16294 2662 16346
rect 2662 16294 2672 16346
rect 2696 16294 2726 16346
rect 2726 16294 2738 16346
rect 2738 16294 2752 16346
rect 2776 16294 2790 16346
rect 2790 16294 2802 16346
rect 2802 16294 2832 16346
rect 2856 16294 2866 16346
rect 2866 16294 2912 16346
rect 2616 16292 2672 16294
rect 2696 16292 2752 16294
rect 2776 16292 2832 16294
rect 2856 16292 2912 16294
rect 7616 16346 7672 16348
rect 7696 16346 7752 16348
rect 7776 16346 7832 16348
rect 7856 16346 7912 16348
rect 7616 16294 7662 16346
rect 7662 16294 7672 16346
rect 7696 16294 7726 16346
rect 7726 16294 7738 16346
rect 7738 16294 7752 16346
rect 7776 16294 7790 16346
rect 7790 16294 7802 16346
rect 7802 16294 7832 16346
rect 7856 16294 7866 16346
rect 7866 16294 7912 16346
rect 7616 16292 7672 16294
rect 7696 16292 7752 16294
rect 7776 16292 7832 16294
rect 7856 16292 7912 16294
rect 12616 16346 12672 16348
rect 12696 16346 12752 16348
rect 12776 16346 12832 16348
rect 12856 16346 12912 16348
rect 12616 16294 12662 16346
rect 12662 16294 12672 16346
rect 12696 16294 12726 16346
rect 12726 16294 12738 16346
rect 12738 16294 12752 16346
rect 12776 16294 12790 16346
rect 12790 16294 12802 16346
rect 12802 16294 12832 16346
rect 12856 16294 12866 16346
rect 12866 16294 12912 16346
rect 12616 16292 12672 16294
rect 12696 16292 12752 16294
rect 12776 16292 12832 16294
rect 12856 16292 12912 16294
rect 17616 16346 17672 16348
rect 17696 16346 17752 16348
rect 17776 16346 17832 16348
rect 17856 16346 17912 16348
rect 17616 16294 17662 16346
rect 17662 16294 17672 16346
rect 17696 16294 17726 16346
rect 17726 16294 17738 16346
rect 17738 16294 17752 16346
rect 17776 16294 17790 16346
rect 17790 16294 17802 16346
rect 17802 16294 17832 16346
rect 17856 16294 17866 16346
rect 17866 16294 17912 16346
rect 17616 16292 17672 16294
rect 17696 16292 17752 16294
rect 17776 16292 17832 16294
rect 17856 16292 17912 16294
rect 22616 16346 22672 16348
rect 22696 16346 22752 16348
rect 22776 16346 22832 16348
rect 22856 16346 22912 16348
rect 22616 16294 22662 16346
rect 22662 16294 22672 16346
rect 22696 16294 22726 16346
rect 22726 16294 22738 16346
rect 22738 16294 22752 16346
rect 22776 16294 22790 16346
rect 22790 16294 22802 16346
rect 22802 16294 22832 16346
rect 22856 16294 22866 16346
rect 22866 16294 22912 16346
rect 22616 16292 22672 16294
rect 22696 16292 22752 16294
rect 22776 16292 22832 16294
rect 22856 16292 22912 16294
rect 27616 16346 27672 16348
rect 27696 16346 27752 16348
rect 27776 16346 27832 16348
rect 27856 16346 27912 16348
rect 27616 16294 27662 16346
rect 27662 16294 27672 16346
rect 27696 16294 27726 16346
rect 27726 16294 27738 16346
rect 27738 16294 27752 16346
rect 27776 16294 27790 16346
rect 27790 16294 27802 16346
rect 27802 16294 27832 16346
rect 27856 16294 27866 16346
rect 27866 16294 27912 16346
rect 27616 16292 27672 16294
rect 27696 16292 27752 16294
rect 27776 16292 27832 16294
rect 27856 16292 27912 16294
rect 32616 16346 32672 16348
rect 32696 16346 32752 16348
rect 32776 16346 32832 16348
rect 32856 16346 32912 16348
rect 32616 16294 32662 16346
rect 32662 16294 32672 16346
rect 32696 16294 32726 16346
rect 32726 16294 32738 16346
rect 32738 16294 32752 16346
rect 32776 16294 32790 16346
rect 32790 16294 32802 16346
rect 32802 16294 32832 16346
rect 32856 16294 32866 16346
rect 32866 16294 32912 16346
rect 32616 16292 32672 16294
rect 32696 16292 32752 16294
rect 32776 16292 32832 16294
rect 32856 16292 32912 16294
rect 37616 16346 37672 16348
rect 37696 16346 37752 16348
rect 37776 16346 37832 16348
rect 37856 16346 37912 16348
rect 37616 16294 37662 16346
rect 37662 16294 37672 16346
rect 37696 16294 37726 16346
rect 37726 16294 37738 16346
rect 37738 16294 37752 16346
rect 37776 16294 37790 16346
rect 37790 16294 37802 16346
rect 37802 16294 37832 16346
rect 37856 16294 37866 16346
rect 37866 16294 37912 16346
rect 37616 16292 37672 16294
rect 37696 16292 37752 16294
rect 37776 16292 37832 16294
rect 37856 16292 37912 16294
rect 1956 15802 2012 15804
rect 2036 15802 2092 15804
rect 2116 15802 2172 15804
rect 2196 15802 2252 15804
rect 1956 15750 2002 15802
rect 2002 15750 2012 15802
rect 2036 15750 2066 15802
rect 2066 15750 2078 15802
rect 2078 15750 2092 15802
rect 2116 15750 2130 15802
rect 2130 15750 2142 15802
rect 2142 15750 2172 15802
rect 2196 15750 2206 15802
rect 2206 15750 2252 15802
rect 1956 15748 2012 15750
rect 2036 15748 2092 15750
rect 2116 15748 2172 15750
rect 2196 15748 2252 15750
rect 6956 15802 7012 15804
rect 7036 15802 7092 15804
rect 7116 15802 7172 15804
rect 7196 15802 7252 15804
rect 6956 15750 7002 15802
rect 7002 15750 7012 15802
rect 7036 15750 7066 15802
rect 7066 15750 7078 15802
rect 7078 15750 7092 15802
rect 7116 15750 7130 15802
rect 7130 15750 7142 15802
rect 7142 15750 7172 15802
rect 7196 15750 7206 15802
rect 7206 15750 7252 15802
rect 6956 15748 7012 15750
rect 7036 15748 7092 15750
rect 7116 15748 7172 15750
rect 7196 15748 7252 15750
rect 11956 15802 12012 15804
rect 12036 15802 12092 15804
rect 12116 15802 12172 15804
rect 12196 15802 12252 15804
rect 11956 15750 12002 15802
rect 12002 15750 12012 15802
rect 12036 15750 12066 15802
rect 12066 15750 12078 15802
rect 12078 15750 12092 15802
rect 12116 15750 12130 15802
rect 12130 15750 12142 15802
rect 12142 15750 12172 15802
rect 12196 15750 12206 15802
rect 12206 15750 12252 15802
rect 11956 15748 12012 15750
rect 12036 15748 12092 15750
rect 12116 15748 12172 15750
rect 12196 15748 12252 15750
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 17002 15802
rect 17002 15750 17012 15802
rect 17036 15750 17066 15802
rect 17066 15750 17078 15802
rect 17078 15750 17092 15802
rect 17116 15750 17130 15802
rect 17130 15750 17142 15802
rect 17142 15750 17172 15802
rect 17196 15750 17206 15802
rect 17206 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 21956 15802 22012 15804
rect 22036 15802 22092 15804
rect 22116 15802 22172 15804
rect 22196 15802 22252 15804
rect 21956 15750 22002 15802
rect 22002 15750 22012 15802
rect 22036 15750 22066 15802
rect 22066 15750 22078 15802
rect 22078 15750 22092 15802
rect 22116 15750 22130 15802
rect 22130 15750 22142 15802
rect 22142 15750 22172 15802
rect 22196 15750 22206 15802
rect 22206 15750 22252 15802
rect 21956 15748 22012 15750
rect 22036 15748 22092 15750
rect 22116 15748 22172 15750
rect 22196 15748 22252 15750
rect 26956 15802 27012 15804
rect 27036 15802 27092 15804
rect 27116 15802 27172 15804
rect 27196 15802 27252 15804
rect 26956 15750 27002 15802
rect 27002 15750 27012 15802
rect 27036 15750 27066 15802
rect 27066 15750 27078 15802
rect 27078 15750 27092 15802
rect 27116 15750 27130 15802
rect 27130 15750 27142 15802
rect 27142 15750 27172 15802
rect 27196 15750 27206 15802
rect 27206 15750 27252 15802
rect 26956 15748 27012 15750
rect 27036 15748 27092 15750
rect 27116 15748 27172 15750
rect 27196 15748 27252 15750
rect 31956 15802 32012 15804
rect 32036 15802 32092 15804
rect 32116 15802 32172 15804
rect 32196 15802 32252 15804
rect 31956 15750 32002 15802
rect 32002 15750 32012 15802
rect 32036 15750 32066 15802
rect 32066 15750 32078 15802
rect 32078 15750 32092 15802
rect 32116 15750 32130 15802
rect 32130 15750 32142 15802
rect 32142 15750 32172 15802
rect 32196 15750 32206 15802
rect 32206 15750 32252 15802
rect 31956 15748 32012 15750
rect 32036 15748 32092 15750
rect 32116 15748 32172 15750
rect 32196 15748 32252 15750
rect 36956 15802 37012 15804
rect 37036 15802 37092 15804
rect 37116 15802 37172 15804
rect 37196 15802 37252 15804
rect 36956 15750 37002 15802
rect 37002 15750 37012 15802
rect 37036 15750 37066 15802
rect 37066 15750 37078 15802
rect 37078 15750 37092 15802
rect 37116 15750 37130 15802
rect 37130 15750 37142 15802
rect 37142 15750 37172 15802
rect 37196 15750 37206 15802
rect 37206 15750 37252 15802
rect 36956 15748 37012 15750
rect 37036 15748 37092 15750
rect 37116 15748 37172 15750
rect 37196 15748 37252 15750
rect 2616 15258 2672 15260
rect 2696 15258 2752 15260
rect 2776 15258 2832 15260
rect 2856 15258 2912 15260
rect 2616 15206 2662 15258
rect 2662 15206 2672 15258
rect 2696 15206 2726 15258
rect 2726 15206 2738 15258
rect 2738 15206 2752 15258
rect 2776 15206 2790 15258
rect 2790 15206 2802 15258
rect 2802 15206 2832 15258
rect 2856 15206 2866 15258
rect 2866 15206 2912 15258
rect 2616 15204 2672 15206
rect 2696 15204 2752 15206
rect 2776 15204 2832 15206
rect 2856 15204 2912 15206
rect 7616 15258 7672 15260
rect 7696 15258 7752 15260
rect 7776 15258 7832 15260
rect 7856 15258 7912 15260
rect 7616 15206 7662 15258
rect 7662 15206 7672 15258
rect 7696 15206 7726 15258
rect 7726 15206 7738 15258
rect 7738 15206 7752 15258
rect 7776 15206 7790 15258
rect 7790 15206 7802 15258
rect 7802 15206 7832 15258
rect 7856 15206 7866 15258
rect 7866 15206 7912 15258
rect 7616 15204 7672 15206
rect 7696 15204 7752 15206
rect 7776 15204 7832 15206
rect 7856 15204 7912 15206
rect 12616 15258 12672 15260
rect 12696 15258 12752 15260
rect 12776 15258 12832 15260
rect 12856 15258 12912 15260
rect 12616 15206 12662 15258
rect 12662 15206 12672 15258
rect 12696 15206 12726 15258
rect 12726 15206 12738 15258
rect 12738 15206 12752 15258
rect 12776 15206 12790 15258
rect 12790 15206 12802 15258
rect 12802 15206 12832 15258
rect 12856 15206 12866 15258
rect 12866 15206 12912 15258
rect 12616 15204 12672 15206
rect 12696 15204 12752 15206
rect 12776 15204 12832 15206
rect 12856 15204 12912 15206
rect 17616 15258 17672 15260
rect 17696 15258 17752 15260
rect 17776 15258 17832 15260
rect 17856 15258 17912 15260
rect 17616 15206 17662 15258
rect 17662 15206 17672 15258
rect 17696 15206 17726 15258
rect 17726 15206 17738 15258
rect 17738 15206 17752 15258
rect 17776 15206 17790 15258
rect 17790 15206 17802 15258
rect 17802 15206 17832 15258
rect 17856 15206 17866 15258
rect 17866 15206 17912 15258
rect 17616 15204 17672 15206
rect 17696 15204 17752 15206
rect 17776 15204 17832 15206
rect 17856 15204 17912 15206
rect 22616 15258 22672 15260
rect 22696 15258 22752 15260
rect 22776 15258 22832 15260
rect 22856 15258 22912 15260
rect 22616 15206 22662 15258
rect 22662 15206 22672 15258
rect 22696 15206 22726 15258
rect 22726 15206 22738 15258
rect 22738 15206 22752 15258
rect 22776 15206 22790 15258
rect 22790 15206 22802 15258
rect 22802 15206 22832 15258
rect 22856 15206 22866 15258
rect 22866 15206 22912 15258
rect 22616 15204 22672 15206
rect 22696 15204 22752 15206
rect 22776 15204 22832 15206
rect 22856 15204 22912 15206
rect 27616 15258 27672 15260
rect 27696 15258 27752 15260
rect 27776 15258 27832 15260
rect 27856 15258 27912 15260
rect 27616 15206 27662 15258
rect 27662 15206 27672 15258
rect 27696 15206 27726 15258
rect 27726 15206 27738 15258
rect 27738 15206 27752 15258
rect 27776 15206 27790 15258
rect 27790 15206 27802 15258
rect 27802 15206 27832 15258
rect 27856 15206 27866 15258
rect 27866 15206 27912 15258
rect 27616 15204 27672 15206
rect 27696 15204 27752 15206
rect 27776 15204 27832 15206
rect 27856 15204 27912 15206
rect 32616 15258 32672 15260
rect 32696 15258 32752 15260
rect 32776 15258 32832 15260
rect 32856 15258 32912 15260
rect 32616 15206 32662 15258
rect 32662 15206 32672 15258
rect 32696 15206 32726 15258
rect 32726 15206 32738 15258
rect 32738 15206 32752 15258
rect 32776 15206 32790 15258
rect 32790 15206 32802 15258
rect 32802 15206 32832 15258
rect 32856 15206 32866 15258
rect 32866 15206 32912 15258
rect 32616 15204 32672 15206
rect 32696 15204 32752 15206
rect 32776 15204 32832 15206
rect 32856 15204 32912 15206
rect 37616 15258 37672 15260
rect 37696 15258 37752 15260
rect 37776 15258 37832 15260
rect 37856 15258 37912 15260
rect 37616 15206 37662 15258
rect 37662 15206 37672 15258
rect 37696 15206 37726 15258
rect 37726 15206 37738 15258
rect 37738 15206 37752 15258
rect 37776 15206 37790 15258
rect 37790 15206 37802 15258
rect 37802 15206 37832 15258
rect 37856 15206 37866 15258
rect 37866 15206 37912 15258
rect 37616 15204 37672 15206
rect 37696 15204 37752 15206
rect 37776 15204 37832 15206
rect 37856 15204 37912 15206
rect 1956 14714 2012 14716
rect 2036 14714 2092 14716
rect 2116 14714 2172 14716
rect 2196 14714 2252 14716
rect 1956 14662 2002 14714
rect 2002 14662 2012 14714
rect 2036 14662 2066 14714
rect 2066 14662 2078 14714
rect 2078 14662 2092 14714
rect 2116 14662 2130 14714
rect 2130 14662 2142 14714
rect 2142 14662 2172 14714
rect 2196 14662 2206 14714
rect 2206 14662 2252 14714
rect 1956 14660 2012 14662
rect 2036 14660 2092 14662
rect 2116 14660 2172 14662
rect 2196 14660 2252 14662
rect 6956 14714 7012 14716
rect 7036 14714 7092 14716
rect 7116 14714 7172 14716
rect 7196 14714 7252 14716
rect 6956 14662 7002 14714
rect 7002 14662 7012 14714
rect 7036 14662 7066 14714
rect 7066 14662 7078 14714
rect 7078 14662 7092 14714
rect 7116 14662 7130 14714
rect 7130 14662 7142 14714
rect 7142 14662 7172 14714
rect 7196 14662 7206 14714
rect 7206 14662 7252 14714
rect 6956 14660 7012 14662
rect 7036 14660 7092 14662
rect 7116 14660 7172 14662
rect 7196 14660 7252 14662
rect 11956 14714 12012 14716
rect 12036 14714 12092 14716
rect 12116 14714 12172 14716
rect 12196 14714 12252 14716
rect 11956 14662 12002 14714
rect 12002 14662 12012 14714
rect 12036 14662 12066 14714
rect 12066 14662 12078 14714
rect 12078 14662 12092 14714
rect 12116 14662 12130 14714
rect 12130 14662 12142 14714
rect 12142 14662 12172 14714
rect 12196 14662 12206 14714
rect 12206 14662 12252 14714
rect 11956 14660 12012 14662
rect 12036 14660 12092 14662
rect 12116 14660 12172 14662
rect 12196 14660 12252 14662
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 17002 14714
rect 17002 14662 17012 14714
rect 17036 14662 17066 14714
rect 17066 14662 17078 14714
rect 17078 14662 17092 14714
rect 17116 14662 17130 14714
rect 17130 14662 17142 14714
rect 17142 14662 17172 14714
rect 17196 14662 17206 14714
rect 17206 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 21956 14714 22012 14716
rect 22036 14714 22092 14716
rect 22116 14714 22172 14716
rect 22196 14714 22252 14716
rect 21956 14662 22002 14714
rect 22002 14662 22012 14714
rect 22036 14662 22066 14714
rect 22066 14662 22078 14714
rect 22078 14662 22092 14714
rect 22116 14662 22130 14714
rect 22130 14662 22142 14714
rect 22142 14662 22172 14714
rect 22196 14662 22206 14714
rect 22206 14662 22252 14714
rect 21956 14660 22012 14662
rect 22036 14660 22092 14662
rect 22116 14660 22172 14662
rect 22196 14660 22252 14662
rect 26956 14714 27012 14716
rect 27036 14714 27092 14716
rect 27116 14714 27172 14716
rect 27196 14714 27252 14716
rect 26956 14662 27002 14714
rect 27002 14662 27012 14714
rect 27036 14662 27066 14714
rect 27066 14662 27078 14714
rect 27078 14662 27092 14714
rect 27116 14662 27130 14714
rect 27130 14662 27142 14714
rect 27142 14662 27172 14714
rect 27196 14662 27206 14714
rect 27206 14662 27252 14714
rect 26956 14660 27012 14662
rect 27036 14660 27092 14662
rect 27116 14660 27172 14662
rect 27196 14660 27252 14662
rect 31956 14714 32012 14716
rect 32036 14714 32092 14716
rect 32116 14714 32172 14716
rect 32196 14714 32252 14716
rect 31956 14662 32002 14714
rect 32002 14662 32012 14714
rect 32036 14662 32066 14714
rect 32066 14662 32078 14714
rect 32078 14662 32092 14714
rect 32116 14662 32130 14714
rect 32130 14662 32142 14714
rect 32142 14662 32172 14714
rect 32196 14662 32206 14714
rect 32206 14662 32252 14714
rect 31956 14660 32012 14662
rect 32036 14660 32092 14662
rect 32116 14660 32172 14662
rect 32196 14660 32252 14662
rect 36956 14714 37012 14716
rect 37036 14714 37092 14716
rect 37116 14714 37172 14716
rect 37196 14714 37252 14716
rect 36956 14662 37002 14714
rect 37002 14662 37012 14714
rect 37036 14662 37066 14714
rect 37066 14662 37078 14714
rect 37078 14662 37092 14714
rect 37116 14662 37130 14714
rect 37130 14662 37142 14714
rect 37142 14662 37172 14714
rect 37196 14662 37206 14714
rect 37206 14662 37252 14714
rect 36956 14660 37012 14662
rect 37036 14660 37092 14662
rect 37116 14660 37172 14662
rect 37196 14660 37252 14662
rect 2616 14170 2672 14172
rect 2696 14170 2752 14172
rect 2776 14170 2832 14172
rect 2856 14170 2912 14172
rect 2616 14118 2662 14170
rect 2662 14118 2672 14170
rect 2696 14118 2726 14170
rect 2726 14118 2738 14170
rect 2738 14118 2752 14170
rect 2776 14118 2790 14170
rect 2790 14118 2802 14170
rect 2802 14118 2832 14170
rect 2856 14118 2866 14170
rect 2866 14118 2912 14170
rect 2616 14116 2672 14118
rect 2696 14116 2752 14118
rect 2776 14116 2832 14118
rect 2856 14116 2912 14118
rect 7616 14170 7672 14172
rect 7696 14170 7752 14172
rect 7776 14170 7832 14172
rect 7856 14170 7912 14172
rect 7616 14118 7662 14170
rect 7662 14118 7672 14170
rect 7696 14118 7726 14170
rect 7726 14118 7738 14170
rect 7738 14118 7752 14170
rect 7776 14118 7790 14170
rect 7790 14118 7802 14170
rect 7802 14118 7832 14170
rect 7856 14118 7866 14170
rect 7866 14118 7912 14170
rect 7616 14116 7672 14118
rect 7696 14116 7752 14118
rect 7776 14116 7832 14118
rect 7856 14116 7912 14118
rect 12616 14170 12672 14172
rect 12696 14170 12752 14172
rect 12776 14170 12832 14172
rect 12856 14170 12912 14172
rect 12616 14118 12662 14170
rect 12662 14118 12672 14170
rect 12696 14118 12726 14170
rect 12726 14118 12738 14170
rect 12738 14118 12752 14170
rect 12776 14118 12790 14170
rect 12790 14118 12802 14170
rect 12802 14118 12832 14170
rect 12856 14118 12866 14170
rect 12866 14118 12912 14170
rect 12616 14116 12672 14118
rect 12696 14116 12752 14118
rect 12776 14116 12832 14118
rect 12856 14116 12912 14118
rect 17616 14170 17672 14172
rect 17696 14170 17752 14172
rect 17776 14170 17832 14172
rect 17856 14170 17912 14172
rect 17616 14118 17662 14170
rect 17662 14118 17672 14170
rect 17696 14118 17726 14170
rect 17726 14118 17738 14170
rect 17738 14118 17752 14170
rect 17776 14118 17790 14170
rect 17790 14118 17802 14170
rect 17802 14118 17832 14170
rect 17856 14118 17866 14170
rect 17866 14118 17912 14170
rect 17616 14116 17672 14118
rect 17696 14116 17752 14118
rect 17776 14116 17832 14118
rect 17856 14116 17912 14118
rect 22616 14170 22672 14172
rect 22696 14170 22752 14172
rect 22776 14170 22832 14172
rect 22856 14170 22912 14172
rect 22616 14118 22662 14170
rect 22662 14118 22672 14170
rect 22696 14118 22726 14170
rect 22726 14118 22738 14170
rect 22738 14118 22752 14170
rect 22776 14118 22790 14170
rect 22790 14118 22802 14170
rect 22802 14118 22832 14170
rect 22856 14118 22866 14170
rect 22866 14118 22912 14170
rect 22616 14116 22672 14118
rect 22696 14116 22752 14118
rect 22776 14116 22832 14118
rect 22856 14116 22912 14118
rect 27616 14170 27672 14172
rect 27696 14170 27752 14172
rect 27776 14170 27832 14172
rect 27856 14170 27912 14172
rect 27616 14118 27662 14170
rect 27662 14118 27672 14170
rect 27696 14118 27726 14170
rect 27726 14118 27738 14170
rect 27738 14118 27752 14170
rect 27776 14118 27790 14170
rect 27790 14118 27802 14170
rect 27802 14118 27832 14170
rect 27856 14118 27866 14170
rect 27866 14118 27912 14170
rect 27616 14116 27672 14118
rect 27696 14116 27752 14118
rect 27776 14116 27832 14118
rect 27856 14116 27912 14118
rect 32616 14170 32672 14172
rect 32696 14170 32752 14172
rect 32776 14170 32832 14172
rect 32856 14170 32912 14172
rect 32616 14118 32662 14170
rect 32662 14118 32672 14170
rect 32696 14118 32726 14170
rect 32726 14118 32738 14170
rect 32738 14118 32752 14170
rect 32776 14118 32790 14170
rect 32790 14118 32802 14170
rect 32802 14118 32832 14170
rect 32856 14118 32866 14170
rect 32866 14118 32912 14170
rect 32616 14116 32672 14118
rect 32696 14116 32752 14118
rect 32776 14116 32832 14118
rect 32856 14116 32912 14118
rect 37616 14170 37672 14172
rect 37696 14170 37752 14172
rect 37776 14170 37832 14172
rect 37856 14170 37912 14172
rect 37616 14118 37662 14170
rect 37662 14118 37672 14170
rect 37696 14118 37726 14170
rect 37726 14118 37738 14170
rect 37738 14118 37752 14170
rect 37776 14118 37790 14170
rect 37790 14118 37802 14170
rect 37802 14118 37832 14170
rect 37856 14118 37866 14170
rect 37866 14118 37912 14170
rect 37616 14116 37672 14118
rect 37696 14116 37752 14118
rect 37776 14116 37832 14118
rect 37856 14116 37912 14118
rect 1956 13626 2012 13628
rect 2036 13626 2092 13628
rect 2116 13626 2172 13628
rect 2196 13626 2252 13628
rect 1956 13574 2002 13626
rect 2002 13574 2012 13626
rect 2036 13574 2066 13626
rect 2066 13574 2078 13626
rect 2078 13574 2092 13626
rect 2116 13574 2130 13626
rect 2130 13574 2142 13626
rect 2142 13574 2172 13626
rect 2196 13574 2206 13626
rect 2206 13574 2252 13626
rect 1956 13572 2012 13574
rect 2036 13572 2092 13574
rect 2116 13572 2172 13574
rect 2196 13572 2252 13574
rect 6956 13626 7012 13628
rect 7036 13626 7092 13628
rect 7116 13626 7172 13628
rect 7196 13626 7252 13628
rect 6956 13574 7002 13626
rect 7002 13574 7012 13626
rect 7036 13574 7066 13626
rect 7066 13574 7078 13626
rect 7078 13574 7092 13626
rect 7116 13574 7130 13626
rect 7130 13574 7142 13626
rect 7142 13574 7172 13626
rect 7196 13574 7206 13626
rect 7206 13574 7252 13626
rect 6956 13572 7012 13574
rect 7036 13572 7092 13574
rect 7116 13572 7172 13574
rect 7196 13572 7252 13574
rect 11956 13626 12012 13628
rect 12036 13626 12092 13628
rect 12116 13626 12172 13628
rect 12196 13626 12252 13628
rect 11956 13574 12002 13626
rect 12002 13574 12012 13626
rect 12036 13574 12066 13626
rect 12066 13574 12078 13626
rect 12078 13574 12092 13626
rect 12116 13574 12130 13626
rect 12130 13574 12142 13626
rect 12142 13574 12172 13626
rect 12196 13574 12206 13626
rect 12206 13574 12252 13626
rect 11956 13572 12012 13574
rect 12036 13572 12092 13574
rect 12116 13572 12172 13574
rect 12196 13572 12252 13574
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 17002 13626
rect 17002 13574 17012 13626
rect 17036 13574 17066 13626
rect 17066 13574 17078 13626
rect 17078 13574 17092 13626
rect 17116 13574 17130 13626
rect 17130 13574 17142 13626
rect 17142 13574 17172 13626
rect 17196 13574 17206 13626
rect 17206 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 21956 13626 22012 13628
rect 22036 13626 22092 13628
rect 22116 13626 22172 13628
rect 22196 13626 22252 13628
rect 21956 13574 22002 13626
rect 22002 13574 22012 13626
rect 22036 13574 22066 13626
rect 22066 13574 22078 13626
rect 22078 13574 22092 13626
rect 22116 13574 22130 13626
rect 22130 13574 22142 13626
rect 22142 13574 22172 13626
rect 22196 13574 22206 13626
rect 22206 13574 22252 13626
rect 21956 13572 22012 13574
rect 22036 13572 22092 13574
rect 22116 13572 22172 13574
rect 22196 13572 22252 13574
rect 26956 13626 27012 13628
rect 27036 13626 27092 13628
rect 27116 13626 27172 13628
rect 27196 13626 27252 13628
rect 26956 13574 27002 13626
rect 27002 13574 27012 13626
rect 27036 13574 27066 13626
rect 27066 13574 27078 13626
rect 27078 13574 27092 13626
rect 27116 13574 27130 13626
rect 27130 13574 27142 13626
rect 27142 13574 27172 13626
rect 27196 13574 27206 13626
rect 27206 13574 27252 13626
rect 26956 13572 27012 13574
rect 27036 13572 27092 13574
rect 27116 13572 27172 13574
rect 27196 13572 27252 13574
rect 31956 13626 32012 13628
rect 32036 13626 32092 13628
rect 32116 13626 32172 13628
rect 32196 13626 32252 13628
rect 31956 13574 32002 13626
rect 32002 13574 32012 13626
rect 32036 13574 32066 13626
rect 32066 13574 32078 13626
rect 32078 13574 32092 13626
rect 32116 13574 32130 13626
rect 32130 13574 32142 13626
rect 32142 13574 32172 13626
rect 32196 13574 32206 13626
rect 32206 13574 32252 13626
rect 31956 13572 32012 13574
rect 32036 13572 32092 13574
rect 32116 13572 32172 13574
rect 32196 13572 32252 13574
rect 36956 13626 37012 13628
rect 37036 13626 37092 13628
rect 37116 13626 37172 13628
rect 37196 13626 37252 13628
rect 36956 13574 37002 13626
rect 37002 13574 37012 13626
rect 37036 13574 37066 13626
rect 37066 13574 37078 13626
rect 37078 13574 37092 13626
rect 37116 13574 37130 13626
rect 37130 13574 37142 13626
rect 37142 13574 37172 13626
rect 37196 13574 37206 13626
rect 37206 13574 37252 13626
rect 36956 13572 37012 13574
rect 37036 13572 37092 13574
rect 37116 13572 37172 13574
rect 37196 13572 37252 13574
rect 2616 13082 2672 13084
rect 2696 13082 2752 13084
rect 2776 13082 2832 13084
rect 2856 13082 2912 13084
rect 2616 13030 2662 13082
rect 2662 13030 2672 13082
rect 2696 13030 2726 13082
rect 2726 13030 2738 13082
rect 2738 13030 2752 13082
rect 2776 13030 2790 13082
rect 2790 13030 2802 13082
rect 2802 13030 2832 13082
rect 2856 13030 2866 13082
rect 2866 13030 2912 13082
rect 2616 13028 2672 13030
rect 2696 13028 2752 13030
rect 2776 13028 2832 13030
rect 2856 13028 2912 13030
rect 7616 13082 7672 13084
rect 7696 13082 7752 13084
rect 7776 13082 7832 13084
rect 7856 13082 7912 13084
rect 7616 13030 7662 13082
rect 7662 13030 7672 13082
rect 7696 13030 7726 13082
rect 7726 13030 7738 13082
rect 7738 13030 7752 13082
rect 7776 13030 7790 13082
rect 7790 13030 7802 13082
rect 7802 13030 7832 13082
rect 7856 13030 7866 13082
rect 7866 13030 7912 13082
rect 7616 13028 7672 13030
rect 7696 13028 7752 13030
rect 7776 13028 7832 13030
rect 7856 13028 7912 13030
rect 12616 13082 12672 13084
rect 12696 13082 12752 13084
rect 12776 13082 12832 13084
rect 12856 13082 12912 13084
rect 12616 13030 12662 13082
rect 12662 13030 12672 13082
rect 12696 13030 12726 13082
rect 12726 13030 12738 13082
rect 12738 13030 12752 13082
rect 12776 13030 12790 13082
rect 12790 13030 12802 13082
rect 12802 13030 12832 13082
rect 12856 13030 12866 13082
rect 12866 13030 12912 13082
rect 12616 13028 12672 13030
rect 12696 13028 12752 13030
rect 12776 13028 12832 13030
rect 12856 13028 12912 13030
rect 17616 13082 17672 13084
rect 17696 13082 17752 13084
rect 17776 13082 17832 13084
rect 17856 13082 17912 13084
rect 17616 13030 17662 13082
rect 17662 13030 17672 13082
rect 17696 13030 17726 13082
rect 17726 13030 17738 13082
rect 17738 13030 17752 13082
rect 17776 13030 17790 13082
rect 17790 13030 17802 13082
rect 17802 13030 17832 13082
rect 17856 13030 17866 13082
rect 17866 13030 17912 13082
rect 17616 13028 17672 13030
rect 17696 13028 17752 13030
rect 17776 13028 17832 13030
rect 17856 13028 17912 13030
rect 22616 13082 22672 13084
rect 22696 13082 22752 13084
rect 22776 13082 22832 13084
rect 22856 13082 22912 13084
rect 22616 13030 22662 13082
rect 22662 13030 22672 13082
rect 22696 13030 22726 13082
rect 22726 13030 22738 13082
rect 22738 13030 22752 13082
rect 22776 13030 22790 13082
rect 22790 13030 22802 13082
rect 22802 13030 22832 13082
rect 22856 13030 22866 13082
rect 22866 13030 22912 13082
rect 22616 13028 22672 13030
rect 22696 13028 22752 13030
rect 22776 13028 22832 13030
rect 22856 13028 22912 13030
rect 27616 13082 27672 13084
rect 27696 13082 27752 13084
rect 27776 13082 27832 13084
rect 27856 13082 27912 13084
rect 27616 13030 27662 13082
rect 27662 13030 27672 13082
rect 27696 13030 27726 13082
rect 27726 13030 27738 13082
rect 27738 13030 27752 13082
rect 27776 13030 27790 13082
rect 27790 13030 27802 13082
rect 27802 13030 27832 13082
rect 27856 13030 27866 13082
rect 27866 13030 27912 13082
rect 27616 13028 27672 13030
rect 27696 13028 27752 13030
rect 27776 13028 27832 13030
rect 27856 13028 27912 13030
rect 32616 13082 32672 13084
rect 32696 13082 32752 13084
rect 32776 13082 32832 13084
rect 32856 13082 32912 13084
rect 32616 13030 32662 13082
rect 32662 13030 32672 13082
rect 32696 13030 32726 13082
rect 32726 13030 32738 13082
rect 32738 13030 32752 13082
rect 32776 13030 32790 13082
rect 32790 13030 32802 13082
rect 32802 13030 32832 13082
rect 32856 13030 32866 13082
rect 32866 13030 32912 13082
rect 32616 13028 32672 13030
rect 32696 13028 32752 13030
rect 32776 13028 32832 13030
rect 32856 13028 32912 13030
rect 37616 13082 37672 13084
rect 37696 13082 37752 13084
rect 37776 13082 37832 13084
rect 37856 13082 37912 13084
rect 37616 13030 37662 13082
rect 37662 13030 37672 13082
rect 37696 13030 37726 13082
rect 37726 13030 37738 13082
rect 37738 13030 37752 13082
rect 37776 13030 37790 13082
rect 37790 13030 37802 13082
rect 37802 13030 37832 13082
rect 37856 13030 37866 13082
rect 37866 13030 37912 13082
rect 37616 13028 37672 13030
rect 37696 13028 37752 13030
rect 37776 13028 37832 13030
rect 37856 13028 37912 13030
rect 1956 12538 2012 12540
rect 2036 12538 2092 12540
rect 2116 12538 2172 12540
rect 2196 12538 2252 12540
rect 1956 12486 2002 12538
rect 2002 12486 2012 12538
rect 2036 12486 2066 12538
rect 2066 12486 2078 12538
rect 2078 12486 2092 12538
rect 2116 12486 2130 12538
rect 2130 12486 2142 12538
rect 2142 12486 2172 12538
rect 2196 12486 2206 12538
rect 2206 12486 2252 12538
rect 1956 12484 2012 12486
rect 2036 12484 2092 12486
rect 2116 12484 2172 12486
rect 2196 12484 2252 12486
rect 6956 12538 7012 12540
rect 7036 12538 7092 12540
rect 7116 12538 7172 12540
rect 7196 12538 7252 12540
rect 6956 12486 7002 12538
rect 7002 12486 7012 12538
rect 7036 12486 7066 12538
rect 7066 12486 7078 12538
rect 7078 12486 7092 12538
rect 7116 12486 7130 12538
rect 7130 12486 7142 12538
rect 7142 12486 7172 12538
rect 7196 12486 7206 12538
rect 7206 12486 7252 12538
rect 6956 12484 7012 12486
rect 7036 12484 7092 12486
rect 7116 12484 7172 12486
rect 7196 12484 7252 12486
rect 11956 12538 12012 12540
rect 12036 12538 12092 12540
rect 12116 12538 12172 12540
rect 12196 12538 12252 12540
rect 11956 12486 12002 12538
rect 12002 12486 12012 12538
rect 12036 12486 12066 12538
rect 12066 12486 12078 12538
rect 12078 12486 12092 12538
rect 12116 12486 12130 12538
rect 12130 12486 12142 12538
rect 12142 12486 12172 12538
rect 12196 12486 12206 12538
rect 12206 12486 12252 12538
rect 11956 12484 12012 12486
rect 12036 12484 12092 12486
rect 12116 12484 12172 12486
rect 12196 12484 12252 12486
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 17002 12538
rect 17002 12486 17012 12538
rect 17036 12486 17066 12538
rect 17066 12486 17078 12538
rect 17078 12486 17092 12538
rect 17116 12486 17130 12538
rect 17130 12486 17142 12538
rect 17142 12486 17172 12538
rect 17196 12486 17206 12538
rect 17206 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 21956 12538 22012 12540
rect 22036 12538 22092 12540
rect 22116 12538 22172 12540
rect 22196 12538 22252 12540
rect 21956 12486 22002 12538
rect 22002 12486 22012 12538
rect 22036 12486 22066 12538
rect 22066 12486 22078 12538
rect 22078 12486 22092 12538
rect 22116 12486 22130 12538
rect 22130 12486 22142 12538
rect 22142 12486 22172 12538
rect 22196 12486 22206 12538
rect 22206 12486 22252 12538
rect 21956 12484 22012 12486
rect 22036 12484 22092 12486
rect 22116 12484 22172 12486
rect 22196 12484 22252 12486
rect 26956 12538 27012 12540
rect 27036 12538 27092 12540
rect 27116 12538 27172 12540
rect 27196 12538 27252 12540
rect 26956 12486 27002 12538
rect 27002 12486 27012 12538
rect 27036 12486 27066 12538
rect 27066 12486 27078 12538
rect 27078 12486 27092 12538
rect 27116 12486 27130 12538
rect 27130 12486 27142 12538
rect 27142 12486 27172 12538
rect 27196 12486 27206 12538
rect 27206 12486 27252 12538
rect 26956 12484 27012 12486
rect 27036 12484 27092 12486
rect 27116 12484 27172 12486
rect 27196 12484 27252 12486
rect 31956 12538 32012 12540
rect 32036 12538 32092 12540
rect 32116 12538 32172 12540
rect 32196 12538 32252 12540
rect 31956 12486 32002 12538
rect 32002 12486 32012 12538
rect 32036 12486 32066 12538
rect 32066 12486 32078 12538
rect 32078 12486 32092 12538
rect 32116 12486 32130 12538
rect 32130 12486 32142 12538
rect 32142 12486 32172 12538
rect 32196 12486 32206 12538
rect 32206 12486 32252 12538
rect 31956 12484 32012 12486
rect 32036 12484 32092 12486
rect 32116 12484 32172 12486
rect 32196 12484 32252 12486
rect 36956 12538 37012 12540
rect 37036 12538 37092 12540
rect 37116 12538 37172 12540
rect 37196 12538 37252 12540
rect 36956 12486 37002 12538
rect 37002 12486 37012 12538
rect 37036 12486 37066 12538
rect 37066 12486 37078 12538
rect 37078 12486 37092 12538
rect 37116 12486 37130 12538
rect 37130 12486 37142 12538
rect 37142 12486 37172 12538
rect 37196 12486 37206 12538
rect 37206 12486 37252 12538
rect 36956 12484 37012 12486
rect 37036 12484 37092 12486
rect 37116 12484 37172 12486
rect 37196 12484 37252 12486
rect 2616 11994 2672 11996
rect 2696 11994 2752 11996
rect 2776 11994 2832 11996
rect 2856 11994 2912 11996
rect 2616 11942 2662 11994
rect 2662 11942 2672 11994
rect 2696 11942 2726 11994
rect 2726 11942 2738 11994
rect 2738 11942 2752 11994
rect 2776 11942 2790 11994
rect 2790 11942 2802 11994
rect 2802 11942 2832 11994
rect 2856 11942 2866 11994
rect 2866 11942 2912 11994
rect 2616 11940 2672 11942
rect 2696 11940 2752 11942
rect 2776 11940 2832 11942
rect 2856 11940 2912 11942
rect 7616 11994 7672 11996
rect 7696 11994 7752 11996
rect 7776 11994 7832 11996
rect 7856 11994 7912 11996
rect 7616 11942 7662 11994
rect 7662 11942 7672 11994
rect 7696 11942 7726 11994
rect 7726 11942 7738 11994
rect 7738 11942 7752 11994
rect 7776 11942 7790 11994
rect 7790 11942 7802 11994
rect 7802 11942 7832 11994
rect 7856 11942 7866 11994
rect 7866 11942 7912 11994
rect 7616 11940 7672 11942
rect 7696 11940 7752 11942
rect 7776 11940 7832 11942
rect 7856 11940 7912 11942
rect 12616 11994 12672 11996
rect 12696 11994 12752 11996
rect 12776 11994 12832 11996
rect 12856 11994 12912 11996
rect 12616 11942 12662 11994
rect 12662 11942 12672 11994
rect 12696 11942 12726 11994
rect 12726 11942 12738 11994
rect 12738 11942 12752 11994
rect 12776 11942 12790 11994
rect 12790 11942 12802 11994
rect 12802 11942 12832 11994
rect 12856 11942 12866 11994
rect 12866 11942 12912 11994
rect 12616 11940 12672 11942
rect 12696 11940 12752 11942
rect 12776 11940 12832 11942
rect 12856 11940 12912 11942
rect 17616 11994 17672 11996
rect 17696 11994 17752 11996
rect 17776 11994 17832 11996
rect 17856 11994 17912 11996
rect 17616 11942 17662 11994
rect 17662 11942 17672 11994
rect 17696 11942 17726 11994
rect 17726 11942 17738 11994
rect 17738 11942 17752 11994
rect 17776 11942 17790 11994
rect 17790 11942 17802 11994
rect 17802 11942 17832 11994
rect 17856 11942 17866 11994
rect 17866 11942 17912 11994
rect 17616 11940 17672 11942
rect 17696 11940 17752 11942
rect 17776 11940 17832 11942
rect 17856 11940 17912 11942
rect 22616 11994 22672 11996
rect 22696 11994 22752 11996
rect 22776 11994 22832 11996
rect 22856 11994 22912 11996
rect 22616 11942 22662 11994
rect 22662 11942 22672 11994
rect 22696 11942 22726 11994
rect 22726 11942 22738 11994
rect 22738 11942 22752 11994
rect 22776 11942 22790 11994
rect 22790 11942 22802 11994
rect 22802 11942 22832 11994
rect 22856 11942 22866 11994
rect 22866 11942 22912 11994
rect 22616 11940 22672 11942
rect 22696 11940 22752 11942
rect 22776 11940 22832 11942
rect 22856 11940 22912 11942
rect 27616 11994 27672 11996
rect 27696 11994 27752 11996
rect 27776 11994 27832 11996
rect 27856 11994 27912 11996
rect 27616 11942 27662 11994
rect 27662 11942 27672 11994
rect 27696 11942 27726 11994
rect 27726 11942 27738 11994
rect 27738 11942 27752 11994
rect 27776 11942 27790 11994
rect 27790 11942 27802 11994
rect 27802 11942 27832 11994
rect 27856 11942 27866 11994
rect 27866 11942 27912 11994
rect 27616 11940 27672 11942
rect 27696 11940 27752 11942
rect 27776 11940 27832 11942
rect 27856 11940 27912 11942
rect 32616 11994 32672 11996
rect 32696 11994 32752 11996
rect 32776 11994 32832 11996
rect 32856 11994 32912 11996
rect 32616 11942 32662 11994
rect 32662 11942 32672 11994
rect 32696 11942 32726 11994
rect 32726 11942 32738 11994
rect 32738 11942 32752 11994
rect 32776 11942 32790 11994
rect 32790 11942 32802 11994
rect 32802 11942 32832 11994
rect 32856 11942 32866 11994
rect 32866 11942 32912 11994
rect 32616 11940 32672 11942
rect 32696 11940 32752 11942
rect 32776 11940 32832 11942
rect 32856 11940 32912 11942
rect 37616 11994 37672 11996
rect 37696 11994 37752 11996
rect 37776 11994 37832 11996
rect 37856 11994 37912 11996
rect 37616 11942 37662 11994
rect 37662 11942 37672 11994
rect 37696 11942 37726 11994
rect 37726 11942 37738 11994
rect 37738 11942 37752 11994
rect 37776 11942 37790 11994
rect 37790 11942 37802 11994
rect 37802 11942 37832 11994
rect 37856 11942 37866 11994
rect 37866 11942 37912 11994
rect 37616 11940 37672 11942
rect 37696 11940 37752 11942
rect 37776 11940 37832 11942
rect 37856 11940 37912 11942
rect 1956 11450 2012 11452
rect 2036 11450 2092 11452
rect 2116 11450 2172 11452
rect 2196 11450 2252 11452
rect 1956 11398 2002 11450
rect 2002 11398 2012 11450
rect 2036 11398 2066 11450
rect 2066 11398 2078 11450
rect 2078 11398 2092 11450
rect 2116 11398 2130 11450
rect 2130 11398 2142 11450
rect 2142 11398 2172 11450
rect 2196 11398 2206 11450
rect 2206 11398 2252 11450
rect 1956 11396 2012 11398
rect 2036 11396 2092 11398
rect 2116 11396 2172 11398
rect 2196 11396 2252 11398
rect 6956 11450 7012 11452
rect 7036 11450 7092 11452
rect 7116 11450 7172 11452
rect 7196 11450 7252 11452
rect 6956 11398 7002 11450
rect 7002 11398 7012 11450
rect 7036 11398 7066 11450
rect 7066 11398 7078 11450
rect 7078 11398 7092 11450
rect 7116 11398 7130 11450
rect 7130 11398 7142 11450
rect 7142 11398 7172 11450
rect 7196 11398 7206 11450
rect 7206 11398 7252 11450
rect 6956 11396 7012 11398
rect 7036 11396 7092 11398
rect 7116 11396 7172 11398
rect 7196 11396 7252 11398
rect 11956 11450 12012 11452
rect 12036 11450 12092 11452
rect 12116 11450 12172 11452
rect 12196 11450 12252 11452
rect 11956 11398 12002 11450
rect 12002 11398 12012 11450
rect 12036 11398 12066 11450
rect 12066 11398 12078 11450
rect 12078 11398 12092 11450
rect 12116 11398 12130 11450
rect 12130 11398 12142 11450
rect 12142 11398 12172 11450
rect 12196 11398 12206 11450
rect 12206 11398 12252 11450
rect 11956 11396 12012 11398
rect 12036 11396 12092 11398
rect 12116 11396 12172 11398
rect 12196 11396 12252 11398
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 17002 11450
rect 17002 11398 17012 11450
rect 17036 11398 17066 11450
rect 17066 11398 17078 11450
rect 17078 11398 17092 11450
rect 17116 11398 17130 11450
rect 17130 11398 17142 11450
rect 17142 11398 17172 11450
rect 17196 11398 17206 11450
rect 17206 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 21956 11450 22012 11452
rect 22036 11450 22092 11452
rect 22116 11450 22172 11452
rect 22196 11450 22252 11452
rect 21956 11398 22002 11450
rect 22002 11398 22012 11450
rect 22036 11398 22066 11450
rect 22066 11398 22078 11450
rect 22078 11398 22092 11450
rect 22116 11398 22130 11450
rect 22130 11398 22142 11450
rect 22142 11398 22172 11450
rect 22196 11398 22206 11450
rect 22206 11398 22252 11450
rect 21956 11396 22012 11398
rect 22036 11396 22092 11398
rect 22116 11396 22172 11398
rect 22196 11396 22252 11398
rect 26956 11450 27012 11452
rect 27036 11450 27092 11452
rect 27116 11450 27172 11452
rect 27196 11450 27252 11452
rect 26956 11398 27002 11450
rect 27002 11398 27012 11450
rect 27036 11398 27066 11450
rect 27066 11398 27078 11450
rect 27078 11398 27092 11450
rect 27116 11398 27130 11450
rect 27130 11398 27142 11450
rect 27142 11398 27172 11450
rect 27196 11398 27206 11450
rect 27206 11398 27252 11450
rect 26956 11396 27012 11398
rect 27036 11396 27092 11398
rect 27116 11396 27172 11398
rect 27196 11396 27252 11398
rect 31956 11450 32012 11452
rect 32036 11450 32092 11452
rect 32116 11450 32172 11452
rect 32196 11450 32252 11452
rect 31956 11398 32002 11450
rect 32002 11398 32012 11450
rect 32036 11398 32066 11450
rect 32066 11398 32078 11450
rect 32078 11398 32092 11450
rect 32116 11398 32130 11450
rect 32130 11398 32142 11450
rect 32142 11398 32172 11450
rect 32196 11398 32206 11450
rect 32206 11398 32252 11450
rect 31956 11396 32012 11398
rect 32036 11396 32092 11398
rect 32116 11396 32172 11398
rect 32196 11396 32252 11398
rect 36956 11450 37012 11452
rect 37036 11450 37092 11452
rect 37116 11450 37172 11452
rect 37196 11450 37252 11452
rect 36956 11398 37002 11450
rect 37002 11398 37012 11450
rect 37036 11398 37066 11450
rect 37066 11398 37078 11450
rect 37078 11398 37092 11450
rect 37116 11398 37130 11450
rect 37130 11398 37142 11450
rect 37142 11398 37172 11450
rect 37196 11398 37206 11450
rect 37206 11398 37252 11450
rect 36956 11396 37012 11398
rect 37036 11396 37092 11398
rect 37116 11396 37172 11398
rect 37196 11396 37252 11398
rect 2616 10906 2672 10908
rect 2696 10906 2752 10908
rect 2776 10906 2832 10908
rect 2856 10906 2912 10908
rect 2616 10854 2662 10906
rect 2662 10854 2672 10906
rect 2696 10854 2726 10906
rect 2726 10854 2738 10906
rect 2738 10854 2752 10906
rect 2776 10854 2790 10906
rect 2790 10854 2802 10906
rect 2802 10854 2832 10906
rect 2856 10854 2866 10906
rect 2866 10854 2912 10906
rect 2616 10852 2672 10854
rect 2696 10852 2752 10854
rect 2776 10852 2832 10854
rect 2856 10852 2912 10854
rect 7616 10906 7672 10908
rect 7696 10906 7752 10908
rect 7776 10906 7832 10908
rect 7856 10906 7912 10908
rect 7616 10854 7662 10906
rect 7662 10854 7672 10906
rect 7696 10854 7726 10906
rect 7726 10854 7738 10906
rect 7738 10854 7752 10906
rect 7776 10854 7790 10906
rect 7790 10854 7802 10906
rect 7802 10854 7832 10906
rect 7856 10854 7866 10906
rect 7866 10854 7912 10906
rect 7616 10852 7672 10854
rect 7696 10852 7752 10854
rect 7776 10852 7832 10854
rect 7856 10852 7912 10854
rect 12616 10906 12672 10908
rect 12696 10906 12752 10908
rect 12776 10906 12832 10908
rect 12856 10906 12912 10908
rect 12616 10854 12662 10906
rect 12662 10854 12672 10906
rect 12696 10854 12726 10906
rect 12726 10854 12738 10906
rect 12738 10854 12752 10906
rect 12776 10854 12790 10906
rect 12790 10854 12802 10906
rect 12802 10854 12832 10906
rect 12856 10854 12866 10906
rect 12866 10854 12912 10906
rect 12616 10852 12672 10854
rect 12696 10852 12752 10854
rect 12776 10852 12832 10854
rect 12856 10852 12912 10854
rect 17616 10906 17672 10908
rect 17696 10906 17752 10908
rect 17776 10906 17832 10908
rect 17856 10906 17912 10908
rect 17616 10854 17662 10906
rect 17662 10854 17672 10906
rect 17696 10854 17726 10906
rect 17726 10854 17738 10906
rect 17738 10854 17752 10906
rect 17776 10854 17790 10906
rect 17790 10854 17802 10906
rect 17802 10854 17832 10906
rect 17856 10854 17866 10906
rect 17866 10854 17912 10906
rect 17616 10852 17672 10854
rect 17696 10852 17752 10854
rect 17776 10852 17832 10854
rect 17856 10852 17912 10854
rect 22616 10906 22672 10908
rect 22696 10906 22752 10908
rect 22776 10906 22832 10908
rect 22856 10906 22912 10908
rect 22616 10854 22662 10906
rect 22662 10854 22672 10906
rect 22696 10854 22726 10906
rect 22726 10854 22738 10906
rect 22738 10854 22752 10906
rect 22776 10854 22790 10906
rect 22790 10854 22802 10906
rect 22802 10854 22832 10906
rect 22856 10854 22866 10906
rect 22866 10854 22912 10906
rect 22616 10852 22672 10854
rect 22696 10852 22752 10854
rect 22776 10852 22832 10854
rect 22856 10852 22912 10854
rect 27616 10906 27672 10908
rect 27696 10906 27752 10908
rect 27776 10906 27832 10908
rect 27856 10906 27912 10908
rect 27616 10854 27662 10906
rect 27662 10854 27672 10906
rect 27696 10854 27726 10906
rect 27726 10854 27738 10906
rect 27738 10854 27752 10906
rect 27776 10854 27790 10906
rect 27790 10854 27802 10906
rect 27802 10854 27832 10906
rect 27856 10854 27866 10906
rect 27866 10854 27912 10906
rect 27616 10852 27672 10854
rect 27696 10852 27752 10854
rect 27776 10852 27832 10854
rect 27856 10852 27912 10854
rect 32616 10906 32672 10908
rect 32696 10906 32752 10908
rect 32776 10906 32832 10908
rect 32856 10906 32912 10908
rect 32616 10854 32662 10906
rect 32662 10854 32672 10906
rect 32696 10854 32726 10906
rect 32726 10854 32738 10906
rect 32738 10854 32752 10906
rect 32776 10854 32790 10906
rect 32790 10854 32802 10906
rect 32802 10854 32832 10906
rect 32856 10854 32866 10906
rect 32866 10854 32912 10906
rect 32616 10852 32672 10854
rect 32696 10852 32752 10854
rect 32776 10852 32832 10854
rect 32856 10852 32912 10854
rect 37616 10906 37672 10908
rect 37696 10906 37752 10908
rect 37776 10906 37832 10908
rect 37856 10906 37912 10908
rect 37616 10854 37662 10906
rect 37662 10854 37672 10906
rect 37696 10854 37726 10906
rect 37726 10854 37738 10906
rect 37738 10854 37752 10906
rect 37776 10854 37790 10906
rect 37790 10854 37802 10906
rect 37802 10854 37832 10906
rect 37856 10854 37866 10906
rect 37866 10854 37912 10906
rect 37616 10852 37672 10854
rect 37696 10852 37752 10854
rect 37776 10852 37832 10854
rect 37856 10852 37912 10854
rect 1956 10362 2012 10364
rect 2036 10362 2092 10364
rect 2116 10362 2172 10364
rect 2196 10362 2252 10364
rect 1956 10310 2002 10362
rect 2002 10310 2012 10362
rect 2036 10310 2066 10362
rect 2066 10310 2078 10362
rect 2078 10310 2092 10362
rect 2116 10310 2130 10362
rect 2130 10310 2142 10362
rect 2142 10310 2172 10362
rect 2196 10310 2206 10362
rect 2206 10310 2252 10362
rect 1956 10308 2012 10310
rect 2036 10308 2092 10310
rect 2116 10308 2172 10310
rect 2196 10308 2252 10310
rect 6956 10362 7012 10364
rect 7036 10362 7092 10364
rect 7116 10362 7172 10364
rect 7196 10362 7252 10364
rect 6956 10310 7002 10362
rect 7002 10310 7012 10362
rect 7036 10310 7066 10362
rect 7066 10310 7078 10362
rect 7078 10310 7092 10362
rect 7116 10310 7130 10362
rect 7130 10310 7142 10362
rect 7142 10310 7172 10362
rect 7196 10310 7206 10362
rect 7206 10310 7252 10362
rect 6956 10308 7012 10310
rect 7036 10308 7092 10310
rect 7116 10308 7172 10310
rect 7196 10308 7252 10310
rect 11956 10362 12012 10364
rect 12036 10362 12092 10364
rect 12116 10362 12172 10364
rect 12196 10362 12252 10364
rect 11956 10310 12002 10362
rect 12002 10310 12012 10362
rect 12036 10310 12066 10362
rect 12066 10310 12078 10362
rect 12078 10310 12092 10362
rect 12116 10310 12130 10362
rect 12130 10310 12142 10362
rect 12142 10310 12172 10362
rect 12196 10310 12206 10362
rect 12206 10310 12252 10362
rect 11956 10308 12012 10310
rect 12036 10308 12092 10310
rect 12116 10308 12172 10310
rect 12196 10308 12252 10310
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 17002 10362
rect 17002 10310 17012 10362
rect 17036 10310 17066 10362
rect 17066 10310 17078 10362
rect 17078 10310 17092 10362
rect 17116 10310 17130 10362
rect 17130 10310 17142 10362
rect 17142 10310 17172 10362
rect 17196 10310 17206 10362
rect 17206 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 21956 10362 22012 10364
rect 22036 10362 22092 10364
rect 22116 10362 22172 10364
rect 22196 10362 22252 10364
rect 21956 10310 22002 10362
rect 22002 10310 22012 10362
rect 22036 10310 22066 10362
rect 22066 10310 22078 10362
rect 22078 10310 22092 10362
rect 22116 10310 22130 10362
rect 22130 10310 22142 10362
rect 22142 10310 22172 10362
rect 22196 10310 22206 10362
rect 22206 10310 22252 10362
rect 21956 10308 22012 10310
rect 22036 10308 22092 10310
rect 22116 10308 22172 10310
rect 22196 10308 22252 10310
rect 26956 10362 27012 10364
rect 27036 10362 27092 10364
rect 27116 10362 27172 10364
rect 27196 10362 27252 10364
rect 26956 10310 27002 10362
rect 27002 10310 27012 10362
rect 27036 10310 27066 10362
rect 27066 10310 27078 10362
rect 27078 10310 27092 10362
rect 27116 10310 27130 10362
rect 27130 10310 27142 10362
rect 27142 10310 27172 10362
rect 27196 10310 27206 10362
rect 27206 10310 27252 10362
rect 26956 10308 27012 10310
rect 27036 10308 27092 10310
rect 27116 10308 27172 10310
rect 27196 10308 27252 10310
rect 31956 10362 32012 10364
rect 32036 10362 32092 10364
rect 32116 10362 32172 10364
rect 32196 10362 32252 10364
rect 31956 10310 32002 10362
rect 32002 10310 32012 10362
rect 32036 10310 32066 10362
rect 32066 10310 32078 10362
rect 32078 10310 32092 10362
rect 32116 10310 32130 10362
rect 32130 10310 32142 10362
rect 32142 10310 32172 10362
rect 32196 10310 32206 10362
rect 32206 10310 32252 10362
rect 31956 10308 32012 10310
rect 32036 10308 32092 10310
rect 32116 10308 32172 10310
rect 32196 10308 32252 10310
rect 36956 10362 37012 10364
rect 37036 10362 37092 10364
rect 37116 10362 37172 10364
rect 37196 10362 37252 10364
rect 36956 10310 37002 10362
rect 37002 10310 37012 10362
rect 37036 10310 37066 10362
rect 37066 10310 37078 10362
rect 37078 10310 37092 10362
rect 37116 10310 37130 10362
rect 37130 10310 37142 10362
rect 37142 10310 37172 10362
rect 37196 10310 37206 10362
rect 37206 10310 37252 10362
rect 36956 10308 37012 10310
rect 37036 10308 37092 10310
rect 37116 10308 37172 10310
rect 37196 10308 37252 10310
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 7616 9818 7672 9820
rect 7696 9818 7752 9820
rect 7776 9818 7832 9820
rect 7856 9818 7912 9820
rect 7616 9766 7662 9818
rect 7662 9766 7672 9818
rect 7696 9766 7726 9818
rect 7726 9766 7738 9818
rect 7738 9766 7752 9818
rect 7776 9766 7790 9818
rect 7790 9766 7802 9818
rect 7802 9766 7832 9818
rect 7856 9766 7866 9818
rect 7866 9766 7912 9818
rect 7616 9764 7672 9766
rect 7696 9764 7752 9766
rect 7776 9764 7832 9766
rect 7856 9764 7912 9766
rect 12616 9818 12672 9820
rect 12696 9818 12752 9820
rect 12776 9818 12832 9820
rect 12856 9818 12912 9820
rect 12616 9766 12662 9818
rect 12662 9766 12672 9818
rect 12696 9766 12726 9818
rect 12726 9766 12738 9818
rect 12738 9766 12752 9818
rect 12776 9766 12790 9818
rect 12790 9766 12802 9818
rect 12802 9766 12832 9818
rect 12856 9766 12866 9818
rect 12866 9766 12912 9818
rect 12616 9764 12672 9766
rect 12696 9764 12752 9766
rect 12776 9764 12832 9766
rect 12856 9764 12912 9766
rect 17616 9818 17672 9820
rect 17696 9818 17752 9820
rect 17776 9818 17832 9820
rect 17856 9818 17912 9820
rect 17616 9766 17662 9818
rect 17662 9766 17672 9818
rect 17696 9766 17726 9818
rect 17726 9766 17738 9818
rect 17738 9766 17752 9818
rect 17776 9766 17790 9818
rect 17790 9766 17802 9818
rect 17802 9766 17832 9818
rect 17856 9766 17866 9818
rect 17866 9766 17912 9818
rect 17616 9764 17672 9766
rect 17696 9764 17752 9766
rect 17776 9764 17832 9766
rect 17856 9764 17912 9766
rect 22616 9818 22672 9820
rect 22696 9818 22752 9820
rect 22776 9818 22832 9820
rect 22856 9818 22912 9820
rect 22616 9766 22662 9818
rect 22662 9766 22672 9818
rect 22696 9766 22726 9818
rect 22726 9766 22738 9818
rect 22738 9766 22752 9818
rect 22776 9766 22790 9818
rect 22790 9766 22802 9818
rect 22802 9766 22832 9818
rect 22856 9766 22866 9818
rect 22866 9766 22912 9818
rect 22616 9764 22672 9766
rect 22696 9764 22752 9766
rect 22776 9764 22832 9766
rect 22856 9764 22912 9766
rect 27616 9818 27672 9820
rect 27696 9818 27752 9820
rect 27776 9818 27832 9820
rect 27856 9818 27912 9820
rect 27616 9766 27662 9818
rect 27662 9766 27672 9818
rect 27696 9766 27726 9818
rect 27726 9766 27738 9818
rect 27738 9766 27752 9818
rect 27776 9766 27790 9818
rect 27790 9766 27802 9818
rect 27802 9766 27832 9818
rect 27856 9766 27866 9818
rect 27866 9766 27912 9818
rect 27616 9764 27672 9766
rect 27696 9764 27752 9766
rect 27776 9764 27832 9766
rect 27856 9764 27912 9766
rect 32616 9818 32672 9820
rect 32696 9818 32752 9820
rect 32776 9818 32832 9820
rect 32856 9818 32912 9820
rect 32616 9766 32662 9818
rect 32662 9766 32672 9818
rect 32696 9766 32726 9818
rect 32726 9766 32738 9818
rect 32738 9766 32752 9818
rect 32776 9766 32790 9818
rect 32790 9766 32802 9818
rect 32802 9766 32832 9818
rect 32856 9766 32866 9818
rect 32866 9766 32912 9818
rect 32616 9764 32672 9766
rect 32696 9764 32752 9766
rect 32776 9764 32832 9766
rect 32856 9764 32912 9766
rect 37616 9818 37672 9820
rect 37696 9818 37752 9820
rect 37776 9818 37832 9820
rect 37856 9818 37912 9820
rect 37616 9766 37662 9818
rect 37662 9766 37672 9818
rect 37696 9766 37726 9818
rect 37726 9766 37738 9818
rect 37738 9766 37752 9818
rect 37776 9766 37790 9818
rect 37790 9766 37802 9818
rect 37802 9766 37832 9818
rect 37856 9766 37866 9818
rect 37866 9766 37912 9818
rect 37616 9764 37672 9766
rect 37696 9764 37752 9766
rect 37776 9764 37832 9766
rect 37856 9764 37912 9766
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 6956 9274 7012 9276
rect 7036 9274 7092 9276
rect 7116 9274 7172 9276
rect 7196 9274 7252 9276
rect 6956 9222 7002 9274
rect 7002 9222 7012 9274
rect 7036 9222 7066 9274
rect 7066 9222 7078 9274
rect 7078 9222 7092 9274
rect 7116 9222 7130 9274
rect 7130 9222 7142 9274
rect 7142 9222 7172 9274
rect 7196 9222 7206 9274
rect 7206 9222 7252 9274
rect 6956 9220 7012 9222
rect 7036 9220 7092 9222
rect 7116 9220 7172 9222
rect 7196 9220 7252 9222
rect 11956 9274 12012 9276
rect 12036 9274 12092 9276
rect 12116 9274 12172 9276
rect 12196 9274 12252 9276
rect 11956 9222 12002 9274
rect 12002 9222 12012 9274
rect 12036 9222 12066 9274
rect 12066 9222 12078 9274
rect 12078 9222 12092 9274
rect 12116 9222 12130 9274
rect 12130 9222 12142 9274
rect 12142 9222 12172 9274
rect 12196 9222 12206 9274
rect 12206 9222 12252 9274
rect 11956 9220 12012 9222
rect 12036 9220 12092 9222
rect 12116 9220 12172 9222
rect 12196 9220 12252 9222
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 17002 9274
rect 17002 9222 17012 9274
rect 17036 9222 17066 9274
rect 17066 9222 17078 9274
rect 17078 9222 17092 9274
rect 17116 9222 17130 9274
rect 17130 9222 17142 9274
rect 17142 9222 17172 9274
rect 17196 9222 17206 9274
rect 17206 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 21956 9274 22012 9276
rect 22036 9274 22092 9276
rect 22116 9274 22172 9276
rect 22196 9274 22252 9276
rect 21956 9222 22002 9274
rect 22002 9222 22012 9274
rect 22036 9222 22066 9274
rect 22066 9222 22078 9274
rect 22078 9222 22092 9274
rect 22116 9222 22130 9274
rect 22130 9222 22142 9274
rect 22142 9222 22172 9274
rect 22196 9222 22206 9274
rect 22206 9222 22252 9274
rect 21956 9220 22012 9222
rect 22036 9220 22092 9222
rect 22116 9220 22172 9222
rect 22196 9220 22252 9222
rect 26956 9274 27012 9276
rect 27036 9274 27092 9276
rect 27116 9274 27172 9276
rect 27196 9274 27252 9276
rect 26956 9222 27002 9274
rect 27002 9222 27012 9274
rect 27036 9222 27066 9274
rect 27066 9222 27078 9274
rect 27078 9222 27092 9274
rect 27116 9222 27130 9274
rect 27130 9222 27142 9274
rect 27142 9222 27172 9274
rect 27196 9222 27206 9274
rect 27206 9222 27252 9274
rect 26956 9220 27012 9222
rect 27036 9220 27092 9222
rect 27116 9220 27172 9222
rect 27196 9220 27252 9222
rect 31956 9274 32012 9276
rect 32036 9274 32092 9276
rect 32116 9274 32172 9276
rect 32196 9274 32252 9276
rect 31956 9222 32002 9274
rect 32002 9222 32012 9274
rect 32036 9222 32066 9274
rect 32066 9222 32078 9274
rect 32078 9222 32092 9274
rect 32116 9222 32130 9274
rect 32130 9222 32142 9274
rect 32142 9222 32172 9274
rect 32196 9222 32206 9274
rect 32206 9222 32252 9274
rect 31956 9220 32012 9222
rect 32036 9220 32092 9222
rect 32116 9220 32172 9222
rect 32196 9220 32252 9222
rect 36956 9274 37012 9276
rect 37036 9274 37092 9276
rect 37116 9274 37172 9276
rect 37196 9274 37252 9276
rect 36956 9222 37002 9274
rect 37002 9222 37012 9274
rect 37036 9222 37066 9274
rect 37066 9222 37078 9274
rect 37078 9222 37092 9274
rect 37116 9222 37130 9274
rect 37130 9222 37142 9274
rect 37142 9222 37172 9274
rect 37196 9222 37206 9274
rect 37206 9222 37252 9274
rect 36956 9220 37012 9222
rect 37036 9220 37092 9222
rect 37116 9220 37172 9222
rect 37196 9220 37252 9222
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 7616 8730 7672 8732
rect 7696 8730 7752 8732
rect 7776 8730 7832 8732
rect 7856 8730 7912 8732
rect 7616 8678 7662 8730
rect 7662 8678 7672 8730
rect 7696 8678 7726 8730
rect 7726 8678 7738 8730
rect 7738 8678 7752 8730
rect 7776 8678 7790 8730
rect 7790 8678 7802 8730
rect 7802 8678 7832 8730
rect 7856 8678 7866 8730
rect 7866 8678 7912 8730
rect 7616 8676 7672 8678
rect 7696 8676 7752 8678
rect 7776 8676 7832 8678
rect 7856 8676 7912 8678
rect 12616 8730 12672 8732
rect 12696 8730 12752 8732
rect 12776 8730 12832 8732
rect 12856 8730 12912 8732
rect 12616 8678 12662 8730
rect 12662 8678 12672 8730
rect 12696 8678 12726 8730
rect 12726 8678 12738 8730
rect 12738 8678 12752 8730
rect 12776 8678 12790 8730
rect 12790 8678 12802 8730
rect 12802 8678 12832 8730
rect 12856 8678 12866 8730
rect 12866 8678 12912 8730
rect 12616 8676 12672 8678
rect 12696 8676 12752 8678
rect 12776 8676 12832 8678
rect 12856 8676 12912 8678
rect 17616 8730 17672 8732
rect 17696 8730 17752 8732
rect 17776 8730 17832 8732
rect 17856 8730 17912 8732
rect 17616 8678 17662 8730
rect 17662 8678 17672 8730
rect 17696 8678 17726 8730
rect 17726 8678 17738 8730
rect 17738 8678 17752 8730
rect 17776 8678 17790 8730
rect 17790 8678 17802 8730
rect 17802 8678 17832 8730
rect 17856 8678 17866 8730
rect 17866 8678 17912 8730
rect 17616 8676 17672 8678
rect 17696 8676 17752 8678
rect 17776 8676 17832 8678
rect 17856 8676 17912 8678
rect 22616 8730 22672 8732
rect 22696 8730 22752 8732
rect 22776 8730 22832 8732
rect 22856 8730 22912 8732
rect 22616 8678 22662 8730
rect 22662 8678 22672 8730
rect 22696 8678 22726 8730
rect 22726 8678 22738 8730
rect 22738 8678 22752 8730
rect 22776 8678 22790 8730
rect 22790 8678 22802 8730
rect 22802 8678 22832 8730
rect 22856 8678 22866 8730
rect 22866 8678 22912 8730
rect 22616 8676 22672 8678
rect 22696 8676 22752 8678
rect 22776 8676 22832 8678
rect 22856 8676 22912 8678
rect 27616 8730 27672 8732
rect 27696 8730 27752 8732
rect 27776 8730 27832 8732
rect 27856 8730 27912 8732
rect 27616 8678 27662 8730
rect 27662 8678 27672 8730
rect 27696 8678 27726 8730
rect 27726 8678 27738 8730
rect 27738 8678 27752 8730
rect 27776 8678 27790 8730
rect 27790 8678 27802 8730
rect 27802 8678 27832 8730
rect 27856 8678 27866 8730
rect 27866 8678 27912 8730
rect 27616 8676 27672 8678
rect 27696 8676 27752 8678
rect 27776 8676 27832 8678
rect 27856 8676 27912 8678
rect 32616 8730 32672 8732
rect 32696 8730 32752 8732
rect 32776 8730 32832 8732
rect 32856 8730 32912 8732
rect 32616 8678 32662 8730
rect 32662 8678 32672 8730
rect 32696 8678 32726 8730
rect 32726 8678 32738 8730
rect 32738 8678 32752 8730
rect 32776 8678 32790 8730
rect 32790 8678 32802 8730
rect 32802 8678 32832 8730
rect 32856 8678 32866 8730
rect 32866 8678 32912 8730
rect 32616 8676 32672 8678
rect 32696 8676 32752 8678
rect 32776 8676 32832 8678
rect 32856 8676 32912 8678
rect 37616 8730 37672 8732
rect 37696 8730 37752 8732
rect 37776 8730 37832 8732
rect 37856 8730 37912 8732
rect 37616 8678 37662 8730
rect 37662 8678 37672 8730
rect 37696 8678 37726 8730
rect 37726 8678 37738 8730
rect 37738 8678 37752 8730
rect 37776 8678 37790 8730
rect 37790 8678 37802 8730
rect 37802 8678 37832 8730
rect 37856 8678 37866 8730
rect 37866 8678 37912 8730
rect 37616 8676 37672 8678
rect 37696 8676 37752 8678
rect 37776 8676 37832 8678
rect 37856 8676 37912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 6956 8186 7012 8188
rect 7036 8186 7092 8188
rect 7116 8186 7172 8188
rect 7196 8186 7252 8188
rect 6956 8134 7002 8186
rect 7002 8134 7012 8186
rect 7036 8134 7066 8186
rect 7066 8134 7078 8186
rect 7078 8134 7092 8186
rect 7116 8134 7130 8186
rect 7130 8134 7142 8186
rect 7142 8134 7172 8186
rect 7196 8134 7206 8186
rect 7206 8134 7252 8186
rect 6956 8132 7012 8134
rect 7036 8132 7092 8134
rect 7116 8132 7172 8134
rect 7196 8132 7252 8134
rect 11956 8186 12012 8188
rect 12036 8186 12092 8188
rect 12116 8186 12172 8188
rect 12196 8186 12252 8188
rect 11956 8134 12002 8186
rect 12002 8134 12012 8186
rect 12036 8134 12066 8186
rect 12066 8134 12078 8186
rect 12078 8134 12092 8186
rect 12116 8134 12130 8186
rect 12130 8134 12142 8186
rect 12142 8134 12172 8186
rect 12196 8134 12206 8186
rect 12206 8134 12252 8186
rect 11956 8132 12012 8134
rect 12036 8132 12092 8134
rect 12116 8132 12172 8134
rect 12196 8132 12252 8134
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 17002 8186
rect 17002 8134 17012 8186
rect 17036 8134 17066 8186
rect 17066 8134 17078 8186
rect 17078 8134 17092 8186
rect 17116 8134 17130 8186
rect 17130 8134 17142 8186
rect 17142 8134 17172 8186
rect 17196 8134 17206 8186
rect 17206 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 21956 8186 22012 8188
rect 22036 8186 22092 8188
rect 22116 8186 22172 8188
rect 22196 8186 22252 8188
rect 21956 8134 22002 8186
rect 22002 8134 22012 8186
rect 22036 8134 22066 8186
rect 22066 8134 22078 8186
rect 22078 8134 22092 8186
rect 22116 8134 22130 8186
rect 22130 8134 22142 8186
rect 22142 8134 22172 8186
rect 22196 8134 22206 8186
rect 22206 8134 22252 8186
rect 21956 8132 22012 8134
rect 22036 8132 22092 8134
rect 22116 8132 22172 8134
rect 22196 8132 22252 8134
rect 26956 8186 27012 8188
rect 27036 8186 27092 8188
rect 27116 8186 27172 8188
rect 27196 8186 27252 8188
rect 26956 8134 27002 8186
rect 27002 8134 27012 8186
rect 27036 8134 27066 8186
rect 27066 8134 27078 8186
rect 27078 8134 27092 8186
rect 27116 8134 27130 8186
rect 27130 8134 27142 8186
rect 27142 8134 27172 8186
rect 27196 8134 27206 8186
rect 27206 8134 27252 8186
rect 26956 8132 27012 8134
rect 27036 8132 27092 8134
rect 27116 8132 27172 8134
rect 27196 8132 27252 8134
rect 31956 8186 32012 8188
rect 32036 8186 32092 8188
rect 32116 8186 32172 8188
rect 32196 8186 32252 8188
rect 31956 8134 32002 8186
rect 32002 8134 32012 8186
rect 32036 8134 32066 8186
rect 32066 8134 32078 8186
rect 32078 8134 32092 8186
rect 32116 8134 32130 8186
rect 32130 8134 32142 8186
rect 32142 8134 32172 8186
rect 32196 8134 32206 8186
rect 32206 8134 32252 8186
rect 31956 8132 32012 8134
rect 32036 8132 32092 8134
rect 32116 8132 32172 8134
rect 32196 8132 32252 8134
rect 36956 8186 37012 8188
rect 37036 8186 37092 8188
rect 37116 8186 37172 8188
rect 37196 8186 37252 8188
rect 36956 8134 37002 8186
rect 37002 8134 37012 8186
rect 37036 8134 37066 8186
rect 37066 8134 37078 8186
rect 37078 8134 37092 8186
rect 37116 8134 37130 8186
rect 37130 8134 37142 8186
rect 37142 8134 37172 8186
rect 37196 8134 37206 8186
rect 37206 8134 37252 8186
rect 36956 8132 37012 8134
rect 37036 8132 37092 8134
rect 37116 8132 37172 8134
rect 37196 8132 37252 8134
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 7616 7642 7672 7644
rect 7696 7642 7752 7644
rect 7776 7642 7832 7644
rect 7856 7642 7912 7644
rect 7616 7590 7662 7642
rect 7662 7590 7672 7642
rect 7696 7590 7726 7642
rect 7726 7590 7738 7642
rect 7738 7590 7752 7642
rect 7776 7590 7790 7642
rect 7790 7590 7802 7642
rect 7802 7590 7832 7642
rect 7856 7590 7866 7642
rect 7866 7590 7912 7642
rect 7616 7588 7672 7590
rect 7696 7588 7752 7590
rect 7776 7588 7832 7590
rect 7856 7588 7912 7590
rect 12616 7642 12672 7644
rect 12696 7642 12752 7644
rect 12776 7642 12832 7644
rect 12856 7642 12912 7644
rect 12616 7590 12662 7642
rect 12662 7590 12672 7642
rect 12696 7590 12726 7642
rect 12726 7590 12738 7642
rect 12738 7590 12752 7642
rect 12776 7590 12790 7642
rect 12790 7590 12802 7642
rect 12802 7590 12832 7642
rect 12856 7590 12866 7642
rect 12866 7590 12912 7642
rect 12616 7588 12672 7590
rect 12696 7588 12752 7590
rect 12776 7588 12832 7590
rect 12856 7588 12912 7590
rect 17616 7642 17672 7644
rect 17696 7642 17752 7644
rect 17776 7642 17832 7644
rect 17856 7642 17912 7644
rect 17616 7590 17662 7642
rect 17662 7590 17672 7642
rect 17696 7590 17726 7642
rect 17726 7590 17738 7642
rect 17738 7590 17752 7642
rect 17776 7590 17790 7642
rect 17790 7590 17802 7642
rect 17802 7590 17832 7642
rect 17856 7590 17866 7642
rect 17866 7590 17912 7642
rect 17616 7588 17672 7590
rect 17696 7588 17752 7590
rect 17776 7588 17832 7590
rect 17856 7588 17912 7590
rect 22616 7642 22672 7644
rect 22696 7642 22752 7644
rect 22776 7642 22832 7644
rect 22856 7642 22912 7644
rect 22616 7590 22662 7642
rect 22662 7590 22672 7642
rect 22696 7590 22726 7642
rect 22726 7590 22738 7642
rect 22738 7590 22752 7642
rect 22776 7590 22790 7642
rect 22790 7590 22802 7642
rect 22802 7590 22832 7642
rect 22856 7590 22866 7642
rect 22866 7590 22912 7642
rect 22616 7588 22672 7590
rect 22696 7588 22752 7590
rect 22776 7588 22832 7590
rect 22856 7588 22912 7590
rect 27616 7642 27672 7644
rect 27696 7642 27752 7644
rect 27776 7642 27832 7644
rect 27856 7642 27912 7644
rect 27616 7590 27662 7642
rect 27662 7590 27672 7642
rect 27696 7590 27726 7642
rect 27726 7590 27738 7642
rect 27738 7590 27752 7642
rect 27776 7590 27790 7642
rect 27790 7590 27802 7642
rect 27802 7590 27832 7642
rect 27856 7590 27866 7642
rect 27866 7590 27912 7642
rect 27616 7588 27672 7590
rect 27696 7588 27752 7590
rect 27776 7588 27832 7590
rect 27856 7588 27912 7590
rect 32616 7642 32672 7644
rect 32696 7642 32752 7644
rect 32776 7642 32832 7644
rect 32856 7642 32912 7644
rect 32616 7590 32662 7642
rect 32662 7590 32672 7642
rect 32696 7590 32726 7642
rect 32726 7590 32738 7642
rect 32738 7590 32752 7642
rect 32776 7590 32790 7642
rect 32790 7590 32802 7642
rect 32802 7590 32832 7642
rect 32856 7590 32866 7642
rect 32866 7590 32912 7642
rect 32616 7588 32672 7590
rect 32696 7588 32752 7590
rect 32776 7588 32832 7590
rect 32856 7588 32912 7590
rect 37616 7642 37672 7644
rect 37696 7642 37752 7644
rect 37776 7642 37832 7644
rect 37856 7642 37912 7644
rect 37616 7590 37662 7642
rect 37662 7590 37672 7642
rect 37696 7590 37726 7642
rect 37726 7590 37738 7642
rect 37738 7590 37752 7642
rect 37776 7590 37790 7642
rect 37790 7590 37802 7642
rect 37802 7590 37832 7642
rect 37856 7590 37866 7642
rect 37866 7590 37912 7642
rect 37616 7588 37672 7590
rect 37696 7588 37752 7590
rect 37776 7588 37832 7590
rect 37856 7588 37912 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 6956 7098 7012 7100
rect 7036 7098 7092 7100
rect 7116 7098 7172 7100
rect 7196 7098 7252 7100
rect 6956 7046 7002 7098
rect 7002 7046 7012 7098
rect 7036 7046 7066 7098
rect 7066 7046 7078 7098
rect 7078 7046 7092 7098
rect 7116 7046 7130 7098
rect 7130 7046 7142 7098
rect 7142 7046 7172 7098
rect 7196 7046 7206 7098
rect 7206 7046 7252 7098
rect 6956 7044 7012 7046
rect 7036 7044 7092 7046
rect 7116 7044 7172 7046
rect 7196 7044 7252 7046
rect 11956 7098 12012 7100
rect 12036 7098 12092 7100
rect 12116 7098 12172 7100
rect 12196 7098 12252 7100
rect 11956 7046 12002 7098
rect 12002 7046 12012 7098
rect 12036 7046 12066 7098
rect 12066 7046 12078 7098
rect 12078 7046 12092 7098
rect 12116 7046 12130 7098
rect 12130 7046 12142 7098
rect 12142 7046 12172 7098
rect 12196 7046 12206 7098
rect 12206 7046 12252 7098
rect 11956 7044 12012 7046
rect 12036 7044 12092 7046
rect 12116 7044 12172 7046
rect 12196 7044 12252 7046
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 17002 7098
rect 17002 7046 17012 7098
rect 17036 7046 17066 7098
rect 17066 7046 17078 7098
rect 17078 7046 17092 7098
rect 17116 7046 17130 7098
rect 17130 7046 17142 7098
rect 17142 7046 17172 7098
rect 17196 7046 17206 7098
rect 17206 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 21956 7098 22012 7100
rect 22036 7098 22092 7100
rect 22116 7098 22172 7100
rect 22196 7098 22252 7100
rect 21956 7046 22002 7098
rect 22002 7046 22012 7098
rect 22036 7046 22066 7098
rect 22066 7046 22078 7098
rect 22078 7046 22092 7098
rect 22116 7046 22130 7098
rect 22130 7046 22142 7098
rect 22142 7046 22172 7098
rect 22196 7046 22206 7098
rect 22206 7046 22252 7098
rect 21956 7044 22012 7046
rect 22036 7044 22092 7046
rect 22116 7044 22172 7046
rect 22196 7044 22252 7046
rect 26956 7098 27012 7100
rect 27036 7098 27092 7100
rect 27116 7098 27172 7100
rect 27196 7098 27252 7100
rect 26956 7046 27002 7098
rect 27002 7046 27012 7098
rect 27036 7046 27066 7098
rect 27066 7046 27078 7098
rect 27078 7046 27092 7098
rect 27116 7046 27130 7098
rect 27130 7046 27142 7098
rect 27142 7046 27172 7098
rect 27196 7046 27206 7098
rect 27206 7046 27252 7098
rect 26956 7044 27012 7046
rect 27036 7044 27092 7046
rect 27116 7044 27172 7046
rect 27196 7044 27252 7046
rect 31956 7098 32012 7100
rect 32036 7098 32092 7100
rect 32116 7098 32172 7100
rect 32196 7098 32252 7100
rect 31956 7046 32002 7098
rect 32002 7046 32012 7098
rect 32036 7046 32066 7098
rect 32066 7046 32078 7098
rect 32078 7046 32092 7098
rect 32116 7046 32130 7098
rect 32130 7046 32142 7098
rect 32142 7046 32172 7098
rect 32196 7046 32206 7098
rect 32206 7046 32252 7098
rect 31956 7044 32012 7046
rect 32036 7044 32092 7046
rect 32116 7044 32172 7046
rect 32196 7044 32252 7046
rect 36956 7098 37012 7100
rect 37036 7098 37092 7100
rect 37116 7098 37172 7100
rect 37196 7098 37252 7100
rect 36956 7046 37002 7098
rect 37002 7046 37012 7098
rect 37036 7046 37066 7098
rect 37066 7046 37078 7098
rect 37078 7046 37092 7098
rect 37116 7046 37130 7098
rect 37130 7046 37142 7098
rect 37142 7046 37172 7098
rect 37196 7046 37206 7098
rect 37206 7046 37252 7098
rect 36956 7044 37012 7046
rect 37036 7044 37092 7046
rect 37116 7044 37172 7046
rect 37196 7044 37252 7046
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 7616 6554 7672 6556
rect 7696 6554 7752 6556
rect 7776 6554 7832 6556
rect 7856 6554 7912 6556
rect 7616 6502 7662 6554
rect 7662 6502 7672 6554
rect 7696 6502 7726 6554
rect 7726 6502 7738 6554
rect 7738 6502 7752 6554
rect 7776 6502 7790 6554
rect 7790 6502 7802 6554
rect 7802 6502 7832 6554
rect 7856 6502 7866 6554
rect 7866 6502 7912 6554
rect 7616 6500 7672 6502
rect 7696 6500 7752 6502
rect 7776 6500 7832 6502
rect 7856 6500 7912 6502
rect 12616 6554 12672 6556
rect 12696 6554 12752 6556
rect 12776 6554 12832 6556
rect 12856 6554 12912 6556
rect 12616 6502 12662 6554
rect 12662 6502 12672 6554
rect 12696 6502 12726 6554
rect 12726 6502 12738 6554
rect 12738 6502 12752 6554
rect 12776 6502 12790 6554
rect 12790 6502 12802 6554
rect 12802 6502 12832 6554
rect 12856 6502 12866 6554
rect 12866 6502 12912 6554
rect 12616 6500 12672 6502
rect 12696 6500 12752 6502
rect 12776 6500 12832 6502
rect 12856 6500 12912 6502
rect 17616 6554 17672 6556
rect 17696 6554 17752 6556
rect 17776 6554 17832 6556
rect 17856 6554 17912 6556
rect 17616 6502 17662 6554
rect 17662 6502 17672 6554
rect 17696 6502 17726 6554
rect 17726 6502 17738 6554
rect 17738 6502 17752 6554
rect 17776 6502 17790 6554
rect 17790 6502 17802 6554
rect 17802 6502 17832 6554
rect 17856 6502 17866 6554
rect 17866 6502 17912 6554
rect 17616 6500 17672 6502
rect 17696 6500 17752 6502
rect 17776 6500 17832 6502
rect 17856 6500 17912 6502
rect 22616 6554 22672 6556
rect 22696 6554 22752 6556
rect 22776 6554 22832 6556
rect 22856 6554 22912 6556
rect 22616 6502 22662 6554
rect 22662 6502 22672 6554
rect 22696 6502 22726 6554
rect 22726 6502 22738 6554
rect 22738 6502 22752 6554
rect 22776 6502 22790 6554
rect 22790 6502 22802 6554
rect 22802 6502 22832 6554
rect 22856 6502 22866 6554
rect 22866 6502 22912 6554
rect 22616 6500 22672 6502
rect 22696 6500 22752 6502
rect 22776 6500 22832 6502
rect 22856 6500 22912 6502
rect 27616 6554 27672 6556
rect 27696 6554 27752 6556
rect 27776 6554 27832 6556
rect 27856 6554 27912 6556
rect 27616 6502 27662 6554
rect 27662 6502 27672 6554
rect 27696 6502 27726 6554
rect 27726 6502 27738 6554
rect 27738 6502 27752 6554
rect 27776 6502 27790 6554
rect 27790 6502 27802 6554
rect 27802 6502 27832 6554
rect 27856 6502 27866 6554
rect 27866 6502 27912 6554
rect 27616 6500 27672 6502
rect 27696 6500 27752 6502
rect 27776 6500 27832 6502
rect 27856 6500 27912 6502
rect 32616 6554 32672 6556
rect 32696 6554 32752 6556
rect 32776 6554 32832 6556
rect 32856 6554 32912 6556
rect 32616 6502 32662 6554
rect 32662 6502 32672 6554
rect 32696 6502 32726 6554
rect 32726 6502 32738 6554
rect 32738 6502 32752 6554
rect 32776 6502 32790 6554
rect 32790 6502 32802 6554
rect 32802 6502 32832 6554
rect 32856 6502 32866 6554
rect 32866 6502 32912 6554
rect 32616 6500 32672 6502
rect 32696 6500 32752 6502
rect 32776 6500 32832 6502
rect 32856 6500 32912 6502
rect 37616 6554 37672 6556
rect 37696 6554 37752 6556
rect 37776 6554 37832 6556
rect 37856 6554 37912 6556
rect 37616 6502 37662 6554
rect 37662 6502 37672 6554
rect 37696 6502 37726 6554
rect 37726 6502 37738 6554
rect 37738 6502 37752 6554
rect 37776 6502 37790 6554
rect 37790 6502 37802 6554
rect 37802 6502 37832 6554
rect 37856 6502 37866 6554
rect 37866 6502 37912 6554
rect 37616 6500 37672 6502
rect 37696 6500 37752 6502
rect 37776 6500 37832 6502
rect 37856 6500 37912 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 6956 6010 7012 6012
rect 7036 6010 7092 6012
rect 7116 6010 7172 6012
rect 7196 6010 7252 6012
rect 6956 5958 7002 6010
rect 7002 5958 7012 6010
rect 7036 5958 7066 6010
rect 7066 5958 7078 6010
rect 7078 5958 7092 6010
rect 7116 5958 7130 6010
rect 7130 5958 7142 6010
rect 7142 5958 7172 6010
rect 7196 5958 7206 6010
rect 7206 5958 7252 6010
rect 6956 5956 7012 5958
rect 7036 5956 7092 5958
rect 7116 5956 7172 5958
rect 7196 5956 7252 5958
rect 11956 6010 12012 6012
rect 12036 6010 12092 6012
rect 12116 6010 12172 6012
rect 12196 6010 12252 6012
rect 11956 5958 12002 6010
rect 12002 5958 12012 6010
rect 12036 5958 12066 6010
rect 12066 5958 12078 6010
rect 12078 5958 12092 6010
rect 12116 5958 12130 6010
rect 12130 5958 12142 6010
rect 12142 5958 12172 6010
rect 12196 5958 12206 6010
rect 12206 5958 12252 6010
rect 11956 5956 12012 5958
rect 12036 5956 12092 5958
rect 12116 5956 12172 5958
rect 12196 5956 12252 5958
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 17002 6010
rect 17002 5958 17012 6010
rect 17036 5958 17066 6010
rect 17066 5958 17078 6010
rect 17078 5958 17092 6010
rect 17116 5958 17130 6010
rect 17130 5958 17142 6010
rect 17142 5958 17172 6010
rect 17196 5958 17206 6010
rect 17206 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 21956 6010 22012 6012
rect 22036 6010 22092 6012
rect 22116 6010 22172 6012
rect 22196 6010 22252 6012
rect 21956 5958 22002 6010
rect 22002 5958 22012 6010
rect 22036 5958 22066 6010
rect 22066 5958 22078 6010
rect 22078 5958 22092 6010
rect 22116 5958 22130 6010
rect 22130 5958 22142 6010
rect 22142 5958 22172 6010
rect 22196 5958 22206 6010
rect 22206 5958 22252 6010
rect 21956 5956 22012 5958
rect 22036 5956 22092 5958
rect 22116 5956 22172 5958
rect 22196 5956 22252 5958
rect 26956 6010 27012 6012
rect 27036 6010 27092 6012
rect 27116 6010 27172 6012
rect 27196 6010 27252 6012
rect 26956 5958 27002 6010
rect 27002 5958 27012 6010
rect 27036 5958 27066 6010
rect 27066 5958 27078 6010
rect 27078 5958 27092 6010
rect 27116 5958 27130 6010
rect 27130 5958 27142 6010
rect 27142 5958 27172 6010
rect 27196 5958 27206 6010
rect 27206 5958 27252 6010
rect 26956 5956 27012 5958
rect 27036 5956 27092 5958
rect 27116 5956 27172 5958
rect 27196 5956 27252 5958
rect 31956 6010 32012 6012
rect 32036 6010 32092 6012
rect 32116 6010 32172 6012
rect 32196 6010 32252 6012
rect 31956 5958 32002 6010
rect 32002 5958 32012 6010
rect 32036 5958 32066 6010
rect 32066 5958 32078 6010
rect 32078 5958 32092 6010
rect 32116 5958 32130 6010
rect 32130 5958 32142 6010
rect 32142 5958 32172 6010
rect 32196 5958 32206 6010
rect 32206 5958 32252 6010
rect 31956 5956 32012 5958
rect 32036 5956 32092 5958
rect 32116 5956 32172 5958
rect 32196 5956 32252 5958
rect 36956 6010 37012 6012
rect 37036 6010 37092 6012
rect 37116 6010 37172 6012
rect 37196 6010 37252 6012
rect 36956 5958 37002 6010
rect 37002 5958 37012 6010
rect 37036 5958 37066 6010
rect 37066 5958 37078 6010
rect 37078 5958 37092 6010
rect 37116 5958 37130 6010
rect 37130 5958 37142 6010
rect 37142 5958 37172 6010
rect 37196 5958 37206 6010
rect 37206 5958 37252 6010
rect 36956 5956 37012 5958
rect 37036 5956 37092 5958
rect 37116 5956 37172 5958
rect 37196 5956 37252 5958
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 7616 5466 7672 5468
rect 7696 5466 7752 5468
rect 7776 5466 7832 5468
rect 7856 5466 7912 5468
rect 7616 5414 7662 5466
rect 7662 5414 7672 5466
rect 7696 5414 7726 5466
rect 7726 5414 7738 5466
rect 7738 5414 7752 5466
rect 7776 5414 7790 5466
rect 7790 5414 7802 5466
rect 7802 5414 7832 5466
rect 7856 5414 7866 5466
rect 7866 5414 7912 5466
rect 7616 5412 7672 5414
rect 7696 5412 7752 5414
rect 7776 5412 7832 5414
rect 7856 5412 7912 5414
rect 12616 5466 12672 5468
rect 12696 5466 12752 5468
rect 12776 5466 12832 5468
rect 12856 5466 12912 5468
rect 12616 5414 12662 5466
rect 12662 5414 12672 5466
rect 12696 5414 12726 5466
rect 12726 5414 12738 5466
rect 12738 5414 12752 5466
rect 12776 5414 12790 5466
rect 12790 5414 12802 5466
rect 12802 5414 12832 5466
rect 12856 5414 12866 5466
rect 12866 5414 12912 5466
rect 12616 5412 12672 5414
rect 12696 5412 12752 5414
rect 12776 5412 12832 5414
rect 12856 5412 12912 5414
rect 17616 5466 17672 5468
rect 17696 5466 17752 5468
rect 17776 5466 17832 5468
rect 17856 5466 17912 5468
rect 17616 5414 17662 5466
rect 17662 5414 17672 5466
rect 17696 5414 17726 5466
rect 17726 5414 17738 5466
rect 17738 5414 17752 5466
rect 17776 5414 17790 5466
rect 17790 5414 17802 5466
rect 17802 5414 17832 5466
rect 17856 5414 17866 5466
rect 17866 5414 17912 5466
rect 17616 5412 17672 5414
rect 17696 5412 17752 5414
rect 17776 5412 17832 5414
rect 17856 5412 17912 5414
rect 22616 5466 22672 5468
rect 22696 5466 22752 5468
rect 22776 5466 22832 5468
rect 22856 5466 22912 5468
rect 22616 5414 22662 5466
rect 22662 5414 22672 5466
rect 22696 5414 22726 5466
rect 22726 5414 22738 5466
rect 22738 5414 22752 5466
rect 22776 5414 22790 5466
rect 22790 5414 22802 5466
rect 22802 5414 22832 5466
rect 22856 5414 22866 5466
rect 22866 5414 22912 5466
rect 22616 5412 22672 5414
rect 22696 5412 22752 5414
rect 22776 5412 22832 5414
rect 22856 5412 22912 5414
rect 27616 5466 27672 5468
rect 27696 5466 27752 5468
rect 27776 5466 27832 5468
rect 27856 5466 27912 5468
rect 27616 5414 27662 5466
rect 27662 5414 27672 5466
rect 27696 5414 27726 5466
rect 27726 5414 27738 5466
rect 27738 5414 27752 5466
rect 27776 5414 27790 5466
rect 27790 5414 27802 5466
rect 27802 5414 27832 5466
rect 27856 5414 27866 5466
rect 27866 5414 27912 5466
rect 27616 5412 27672 5414
rect 27696 5412 27752 5414
rect 27776 5412 27832 5414
rect 27856 5412 27912 5414
rect 32616 5466 32672 5468
rect 32696 5466 32752 5468
rect 32776 5466 32832 5468
rect 32856 5466 32912 5468
rect 32616 5414 32662 5466
rect 32662 5414 32672 5466
rect 32696 5414 32726 5466
rect 32726 5414 32738 5466
rect 32738 5414 32752 5466
rect 32776 5414 32790 5466
rect 32790 5414 32802 5466
rect 32802 5414 32832 5466
rect 32856 5414 32866 5466
rect 32866 5414 32912 5466
rect 32616 5412 32672 5414
rect 32696 5412 32752 5414
rect 32776 5412 32832 5414
rect 32856 5412 32912 5414
rect 37616 5466 37672 5468
rect 37696 5466 37752 5468
rect 37776 5466 37832 5468
rect 37856 5466 37912 5468
rect 37616 5414 37662 5466
rect 37662 5414 37672 5466
rect 37696 5414 37726 5466
rect 37726 5414 37738 5466
rect 37738 5414 37752 5466
rect 37776 5414 37790 5466
rect 37790 5414 37802 5466
rect 37802 5414 37832 5466
rect 37856 5414 37866 5466
rect 37866 5414 37912 5466
rect 37616 5412 37672 5414
rect 37696 5412 37752 5414
rect 37776 5412 37832 5414
rect 37856 5412 37912 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 6956 4922 7012 4924
rect 7036 4922 7092 4924
rect 7116 4922 7172 4924
rect 7196 4922 7252 4924
rect 6956 4870 7002 4922
rect 7002 4870 7012 4922
rect 7036 4870 7066 4922
rect 7066 4870 7078 4922
rect 7078 4870 7092 4922
rect 7116 4870 7130 4922
rect 7130 4870 7142 4922
rect 7142 4870 7172 4922
rect 7196 4870 7206 4922
rect 7206 4870 7252 4922
rect 6956 4868 7012 4870
rect 7036 4868 7092 4870
rect 7116 4868 7172 4870
rect 7196 4868 7252 4870
rect 11956 4922 12012 4924
rect 12036 4922 12092 4924
rect 12116 4922 12172 4924
rect 12196 4922 12252 4924
rect 11956 4870 12002 4922
rect 12002 4870 12012 4922
rect 12036 4870 12066 4922
rect 12066 4870 12078 4922
rect 12078 4870 12092 4922
rect 12116 4870 12130 4922
rect 12130 4870 12142 4922
rect 12142 4870 12172 4922
rect 12196 4870 12206 4922
rect 12206 4870 12252 4922
rect 11956 4868 12012 4870
rect 12036 4868 12092 4870
rect 12116 4868 12172 4870
rect 12196 4868 12252 4870
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 17002 4922
rect 17002 4870 17012 4922
rect 17036 4870 17066 4922
rect 17066 4870 17078 4922
rect 17078 4870 17092 4922
rect 17116 4870 17130 4922
rect 17130 4870 17142 4922
rect 17142 4870 17172 4922
rect 17196 4870 17206 4922
rect 17206 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 21956 4922 22012 4924
rect 22036 4922 22092 4924
rect 22116 4922 22172 4924
rect 22196 4922 22252 4924
rect 21956 4870 22002 4922
rect 22002 4870 22012 4922
rect 22036 4870 22066 4922
rect 22066 4870 22078 4922
rect 22078 4870 22092 4922
rect 22116 4870 22130 4922
rect 22130 4870 22142 4922
rect 22142 4870 22172 4922
rect 22196 4870 22206 4922
rect 22206 4870 22252 4922
rect 21956 4868 22012 4870
rect 22036 4868 22092 4870
rect 22116 4868 22172 4870
rect 22196 4868 22252 4870
rect 26956 4922 27012 4924
rect 27036 4922 27092 4924
rect 27116 4922 27172 4924
rect 27196 4922 27252 4924
rect 26956 4870 27002 4922
rect 27002 4870 27012 4922
rect 27036 4870 27066 4922
rect 27066 4870 27078 4922
rect 27078 4870 27092 4922
rect 27116 4870 27130 4922
rect 27130 4870 27142 4922
rect 27142 4870 27172 4922
rect 27196 4870 27206 4922
rect 27206 4870 27252 4922
rect 26956 4868 27012 4870
rect 27036 4868 27092 4870
rect 27116 4868 27172 4870
rect 27196 4868 27252 4870
rect 31956 4922 32012 4924
rect 32036 4922 32092 4924
rect 32116 4922 32172 4924
rect 32196 4922 32252 4924
rect 31956 4870 32002 4922
rect 32002 4870 32012 4922
rect 32036 4870 32066 4922
rect 32066 4870 32078 4922
rect 32078 4870 32092 4922
rect 32116 4870 32130 4922
rect 32130 4870 32142 4922
rect 32142 4870 32172 4922
rect 32196 4870 32206 4922
rect 32206 4870 32252 4922
rect 31956 4868 32012 4870
rect 32036 4868 32092 4870
rect 32116 4868 32172 4870
rect 32196 4868 32252 4870
rect 36956 4922 37012 4924
rect 37036 4922 37092 4924
rect 37116 4922 37172 4924
rect 37196 4922 37252 4924
rect 36956 4870 37002 4922
rect 37002 4870 37012 4922
rect 37036 4870 37066 4922
rect 37066 4870 37078 4922
rect 37078 4870 37092 4922
rect 37116 4870 37130 4922
rect 37130 4870 37142 4922
rect 37142 4870 37172 4922
rect 37196 4870 37206 4922
rect 37206 4870 37252 4922
rect 36956 4868 37012 4870
rect 37036 4868 37092 4870
rect 37116 4868 37172 4870
rect 37196 4868 37252 4870
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 7616 4378 7672 4380
rect 7696 4378 7752 4380
rect 7776 4378 7832 4380
rect 7856 4378 7912 4380
rect 7616 4326 7662 4378
rect 7662 4326 7672 4378
rect 7696 4326 7726 4378
rect 7726 4326 7738 4378
rect 7738 4326 7752 4378
rect 7776 4326 7790 4378
rect 7790 4326 7802 4378
rect 7802 4326 7832 4378
rect 7856 4326 7866 4378
rect 7866 4326 7912 4378
rect 7616 4324 7672 4326
rect 7696 4324 7752 4326
rect 7776 4324 7832 4326
rect 7856 4324 7912 4326
rect 12616 4378 12672 4380
rect 12696 4378 12752 4380
rect 12776 4378 12832 4380
rect 12856 4378 12912 4380
rect 12616 4326 12662 4378
rect 12662 4326 12672 4378
rect 12696 4326 12726 4378
rect 12726 4326 12738 4378
rect 12738 4326 12752 4378
rect 12776 4326 12790 4378
rect 12790 4326 12802 4378
rect 12802 4326 12832 4378
rect 12856 4326 12866 4378
rect 12866 4326 12912 4378
rect 12616 4324 12672 4326
rect 12696 4324 12752 4326
rect 12776 4324 12832 4326
rect 12856 4324 12912 4326
rect 17616 4378 17672 4380
rect 17696 4378 17752 4380
rect 17776 4378 17832 4380
rect 17856 4378 17912 4380
rect 17616 4326 17662 4378
rect 17662 4326 17672 4378
rect 17696 4326 17726 4378
rect 17726 4326 17738 4378
rect 17738 4326 17752 4378
rect 17776 4326 17790 4378
rect 17790 4326 17802 4378
rect 17802 4326 17832 4378
rect 17856 4326 17866 4378
rect 17866 4326 17912 4378
rect 17616 4324 17672 4326
rect 17696 4324 17752 4326
rect 17776 4324 17832 4326
rect 17856 4324 17912 4326
rect 22616 4378 22672 4380
rect 22696 4378 22752 4380
rect 22776 4378 22832 4380
rect 22856 4378 22912 4380
rect 22616 4326 22662 4378
rect 22662 4326 22672 4378
rect 22696 4326 22726 4378
rect 22726 4326 22738 4378
rect 22738 4326 22752 4378
rect 22776 4326 22790 4378
rect 22790 4326 22802 4378
rect 22802 4326 22832 4378
rect 22856 4326 22866 4378
rect 22866 4326 22912 4378
rect 22616 4324 22672 4326
rect 22696 4324 22752 4326
rect 22776 4324 22832 4326
rect 22856 4324 22912 4326
rect 27616 4378 27672 4380
rect 27696 4378 27752 4380
rect 27776 4378 27832 4380
rect 27856 4378 27912 4380
rect 27616 4326 27662 4378
rect 27662 4326 27672 4378
rect 27696 4326 27726 4378
rect 27726 4326 27738 4378
rect 27738 4326 27752 4378
rect 27776 4326 27790 4378
rect 27790 4326 27802 4378
rect 27802 4326 27832 4378
rect 27856 4326 27866 4378
rect 27866 4326 27912 4378
rect 27616 4324 27672 4326
rect 27696 4324 27752 4326
rect 27776 4324 27832 4326
rect 27856 4324 27912 4326
rect 32616 4378 32672 4380
rect 32696 4378 32752 4380
rect 32776 4378 32832 4380
rect 32856 4378 32912 4380
rect 32616 4326 32662 4378
rect 32662 4326 32672 4378
rect 32696 4326 32726 4378
rect 32726 4326 32738 4378
rect 32738 4326 32752 4378
rect 32776 4326 32790 4378
rect 32790 4326 32802 4378
rect 32802 4326 32832 4378
rect 32856 4326 32866 4378
rect 32866 4326 32912 4378
rect 32616 4324 32672 4326
rect 32696 4324 32752 4326
rect 32776 4324 32832 4326
rect 32856 4324 32912 4326
rect 37616 4378 37672 4380
rect 37696 4378 37752 4380
rect 37776 4378 37832 4380
rect 37856 4378 37912 4380
rect 37616 4326 37662 4378
rect 37662 4326 37672 4378
rect 37696 4326 37726 4378
rect 37726 4326 37738 4378
rect 37738 4326 37752 4378
rect 37776 4326 37790 4378
rect 37790 4326 37802 4378
rect 37802 4326 37832 4378
rect 37856 4326 37866 4378
rect 37866 4326 37912 4378
rect 37616 4324 37672 4326
rect 37696 4324 37752 4326
rect 37776 4324 37832 4326
rect 37856 4324 37912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 6956 3834 7012 3836
rect 7036 3834 7092 3836
rect 7116 3834 7172 3836
rect 7196 3834 7252 3836
rect 6956 3782 7002 3834
rect 7002 3782 7012 3834
rect 7036 3782 7066 3834
rect 7066 3782 7078 3834
rect 7078 3782 7092 3834
rect 7116 3782 7130 3834
rect 7130 3782 7142 3834
rect 7142 3782 7172 3834
rect 7196 3782 7206 3834
rect 7206 3782 7252 3834
rect 6956 3780 7012 3782
rect 7036 3780 7092 3782
rect 7116 3780 7172 3782
rect 7196 3780 7252 3782
rect 11956 3834 12012 3836
rect 12036 3834 12092 3836
rect 12116 3834 12172 3836
rect 12196 3834 12252 3836
rect 11956 3782 12002 3834
rect 12002 3782 12012 3834
rect 12036 3782 12066 3834
rect 12066 3782 12078 3834
rect 12078 3782 12092 3834
rect 12116 3782 12130 3834
rect 12130 3782 12142 3834
rect 12142 3782 12172 3834
rect 12196 3782 12206 3834
rect 12206 3782 12252 3834
rect 11956 3780 12012 3782
rect 12036 3780 12092 3782
rect 12116 3780 12172 3782
rect 12196 3780 12252 3782
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 17002 3834
rect 17002 3782 17012 3834
rect 17036 3782 17066 3834
rect 17066 3782 17078 3834
rect 17078 3782 17092 3834
rect 17116 3782 17130 3834
rect 17130 3782 17142 3834
rect 17142 3782 17172 3834
rect 17196 3782 17206 3834
rect 17206 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 21956 3834 22012 3836
rect 22036 3834 22092 3836
rect 22116 3834 22172 3836
rect 22196 3834 22252 3836
rect 21956 3782 22002 3834
rect 22002 3782 22012 3834
rect 22036 3782 22066 3834
rect 22066 3782 22078 3834
rect 22078 3782 22092 3834
rect 22116 3782 22130 3834
rect 22130 3782 22142 3834
rect 22142 3782 22172 3834
rect 22196 3782 22206 3834
rect 22206 3782 22252 3834
rect 21956 3780 22012 3782
rect 22036 3780 22092 3782
rect 22116 3780 22172 3782
rect 22196 3780 22252 3782
rect 26956 3834 27012 3836
rect 27036 3834 27092 3836
rect 27116 3834 27172 3836
rect 27196 3834 27252 3836
rect 26956 3782 27002 3834
rect 27002 3782 27012 3834
rect 27036 3782 27066 3834
rect 27066 3782 27078 3834
rect 27078 3782 27092 3834
rect 27116 3782 27130 3834
rect 27130 3782 27142 3834
rect 27142 3782 27172 3834
rect 27196 3782 27206 3834
rect 27206 3782 27252 3834
rect 26956 3780 27012 3782
rect 27036 3780 27092 3782
rect 27116 3780 27172 3782
rect 27196 3780 27252 3782
rect 31956 3834 32012 3836
rect 32036 3834 32092 3836
rect 32116 3834 32172 3836
rect 32196 3834 32252 3836
rect 31956 3782 32002 3834
rect 32002 3782 32012 3834
rect 32036 3782 32066 3834
rect 32066 3782 32078 3834
rect 32078 3782 32092 3834
rect 32116 3782 32130 3834
rect 32130 3782 32142 3834
rect 32142 3782 32172 3834
rect 32196 3782 32206 3834
rect 32206 3782 32252 3834
rect 31956 3780 32012 3782
rect 32036 3780 32092 3782
rect 32116 3780 32172 3782
rect 32196 3780 32252 3782
rect 36956 3834 37012 3836
rect 37036 3834 37092 3836
rect 37116 3834 37172 3836
rect 37196 3834 37252 3836
rect 36956 3782 37002 3834
rect 37002 3782 37012 3834
rect 37036 3782 37066 3834
rect 37066 3782 37078 3834
rect 37078 3782 37092 3834
rect 37116 3782 37130 3834
rect 37130 3782 37142 3834
rect 37142 3782 37172 3834
rect 37196 3782 37206 3834
rect 37206 3782 37252 3834
rect 36956 3780 37012 3782
rect 37036 3780 37092 3782
rect 37116 3780 37172 3782
rect 37196 3780 37252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 7616 3290 7672 3292
rect 7696 3290 7752 3292
rect 7776 3290 7832 3292
rect 7856 3290 7912 3292
rect 7616 3238 7662 3290
rect 7662 3238 7672 3290
rect 7696 3238 7726 3290
rect 7726 3238 7738 3290
rect 7738 3238 7752 3290
rect 7776 3238 7790 3290
rect 7790 3238 7802 3290
rect 7802 3238 7832 3290
rect 7856 3238 7866 3290
rect 7866 3238 7912 3290
rect 7616 3236 7672 3238
rect 7696 3236 7752 3238
rect 7776 3236 7832 3238
rect 7856 3236 7912 3238
rect 12616 3290 12672 3292
rect 12696 3290 12752 3292
rect 12776 3290 12832 3292
rect 12856 3290 12912 3292
rect 12616 3238 12662 3290
rect 12662 3238 12672 3290
rect 12696 3238 12726 3290
rect 12726 3238 12738 3290
rect 12738 3238 12752 3290
rect 12776 3238 12790 3290
rect 12790 3238 12802 3290
rect 12802 3238 12832 3290
rect 12856 3238 12866 3290
rect 12866 3238 12912 3290
rect 12616 3236 12672 3238
rect 12696 3236 12752 3238
rect 12776 3236 12832 3238
rect 12856 3236 12912 3238
rect 17616 3290 17672 3292
rect 17696 3290 17752 3292
rect 17776 3290 17832 3292
rect 17856 3290 17912 3292
rect 17616 3238 17662 3290
rect 17662 3238 17672 3290
rect 17696 3238 17726 3290
rect 17726 3238 17738 3290
rect 17738 3238 17752 3290
rect 17776 3238 17790 3290
rect 17790 3238 17802 3290
rect 17802 3238 17832 3290
rect 17856 3238 17866 3290
rect 17866 3238 17912 3290
rect 17616 3236 17672 3238
rect 17696 3236 17752 3238
rect 17776 3236 17832 3238
rect 17856 3236 17912 3238
rect 22616 3290 22672 3292
rect 22696 3290 22752 3292
rect 22776 3290 22832 3292
rect 22856 3290 22912 3292
rect 22616 3238 22662 3290
rect 22662 3238 22672 3290
rect 22696 3238 22726 3290
rect 22726 3238 22738 3290
rect 22738 3238 22752 3290
rect 22776 3238 22790 3290
rect 22790 3238 22802 3290
rect 22802 3238 22832 3290
rect 22856 3238 22866 3290
rect 22866 3238 22912 3290
rect 22616 3236 22672 3238
rect 22696 3236 22752 3238
rect 22776 3236 22832 3238
rect 22856 3236 22912 3238
rect 27616 3290 27672 3292
rect 27696 3290 27752 3292
rect 27776 3290 27832 3292
rect 27856 3290 27912 3292
rect 27616 3238 27662 3290
rect 27662 3238 27672 3290
rect 27696 3238 27726 3290
rect 27726 3238 27738 3290
rect 27738 3238 27752 3290
rect 27776 3238 27790 3290
rect 27790 3238 27802 3290
rect 27802 3238 27832 3290
rect 27856 3238 27866 3290
rect 27866 3238 27912 3290
rect 27616 3236 27672 3238
rect 27696 3236 27752 3238
rect 27776 3236 27832 3238
rect 27856 3236 27912 3238
rect 32616 3290 32672 3292
rect 32696 3290 32752 3292
rect 32776 3290 32832 3292
rect 32856 3290 32912 3292
rect 32616 3238 32662 3290
rect 32662 3238 32672 3290
rect 32696 3238 32726 3290
rect 32726 3238 32738 3290
rect 32738 3238 32752 3290
rect 32776 3238 32790 3290
rect 32790 3238 32802 3290
rect 32802 3238 32832 3290
rect 32856 3238 32866 3290
rect 32866 3238 32912 3290
rect 32616 3236 32672 3238
rect 32696 3236 32752 3238
rect 32776 3236 32832 3238
rect 32856 3236 32912 3238
rect 37616 3290 37672 3292
rect 37696 3290 37752 3292
rect 37776 3290 37832 3292
rect 37856 3290 37912 3292
rect 37616 3238 37662 3290
rect 37662 3238 37672 3290
rect 37696 3238 37726 3290
rect 37726 3238 37738 3290
rect 37738 3238 37752 3290
rect 37776 3238 37790 3290
rect 37790 3238 37802 3290
rect 37802 3238 37832 3290
rect 37856 3238 37866 3290
rect 37866 3238 37912 3290
rect 37616 3236 37672 3238
rect 37696 3236 37752 3238
rect 37776 3236 37832 3238
rect 37856 3236 37912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 6956 2746 7012 2748
rect 7036 2746 7092 2748
rect 7116 2746 7172 2748
rect 7196 2746 7252 2748
rect 6956 2694 7002 2746
rect 7002 2694 7012 2746
rect 7036 2694 7066 2746
rect 7066 2694 7078 2746
rect 7078 2694 7092 2746
rect 7116 2694 7130 2746
rect 7130 2694 7142 2746
rect 7142 2694 7172 2746
rect 7196 2694 7206 2746
rect 7206 2694 7252 2746
rect 6956 2692 7012 2694
rect 7036 2692 7092 2694
rect 7116 2692 7172 2694
rect 7196 2692 7252 2694
rect 11956 2746 12012 2748
rect 12036 2746 12092 2748
rect 12116 2746 12172 2748
rect 12196 2746 12252 2748
rect 11956 2694 12002 2746
rect 12002 2694 12012 2746
rect 12036 2694 12066 2746
rect 12066 2694 12078 2746
rect 12078 2694 12092 2746
rect 12116 2694 12130 2746
rect 12130 2694 12142 2746
rect 12142 2694 12172 2746
rect 12196 2694 12206 2746
rect 12206 2694 12252 2746
rect 11956 2692 12012 2694
rect 12036 2692 12092 2694
rect 12116 2692 12172 2694
rect 12196 2692 12252 2694
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 17002 2746
rect 17002 2694 17012 2746
rect 17036 2694 17066 2746
rect 17066 2694 17078 2746
rect 17078 2694 17092 2746
rect 17116 2694 17130 2746
rect 17130 2694 17142 2746
rect 17142 2694 17172 2746
rect 17196 2694 17206 2746
rect 17206 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 21956 2746 22012 2748
rect 22036 2746 22092 2748
rect 22116 2746 22172 2748
rect 22196 2746 22252 2748
rect 21956 2694 22002 2746
rect 22002 2694 22012 2746
rect 22036 2694 22066 2746
rect 22066 2694 22078 2746
rect 22078 2694 22092 2746
rect 22116 2694 22130 2746
rect 22130 2694 22142 2746
rect 22142 2694 22172 2746
rect 22196 2694 22206 2746
rect 22206 2694 22252 2746
rect 21956 2692 22012 2694
rect 22036 2692 22092 2694
rect 22116 2692 22172 2694
rect 22196 2692 22252 2694
rect 26956 2746 27012 2748
rect 27036 2746 27092 2748
rect 27116 2746 27172 2748
rect 27196 2746 27252 2748
rect 26956 2694 27002 2746
rect 27002 2694 27012 2746
rect 27036 2694 27066 2746
rect 27066 2694 27078 2746
rect 27078 2694 27092 2746
rect 27116 2694 27130 2746
rect 27130 2694 27142 2746
rect 27142 2694 27172 2746
rect 27196 2694 27206 2746
rect 27206 2694 27252 2746
rect 26956 2692 27012 2694
rect 27036 2692 27092 2694
rect 27116 2692 27172 2694
rect 27196 2692 27252 2694
rect 31956 2746 32012 2748
rect 32036 2746 32092 2748
rect 32116 2746 32172 2748
rect 32196 2746 32252 2748
rect 31956 2694 32002 2746
rect 32002 2694 32012 2746
rect 32036 2694 32066 2746
rect 32066 2694 32078 2746
rect 32078 2694 32092 2746
rect 32116 2694 32130 2746
rect 32130 2694 32142 2746
rect 32142 2694 32172 2746
rect 32196 2694 32206 2746
rect 32206 2694 32252 2746
rect 31956 2692 32012 2694
rect 32036 2692 32092 2694
rect 32116 2692 32172 2694
rect 32196 2692 32252 2694
rect 36956 2746 37012 2748
rect 37036 2746 37092 2748
rect 37116 2746 37172 2748
rect 37196 2746 37252 2748
rect 36956 2694 37002 2746
rect 37002 2694 37012 2746
rect 37036 2694 37066 2746
rect 37066 2694 37078 2746
rect 37078 2694 37092 2746
rect 37116 2694 37130 2746
rect 37130 2694 37142 2746
rect 37142 2694 37172 2746
rect 37196 2694 37206 2746
rect 37206 2694 37252 2746
rect 36956 2692 37012 2694
rect 37036 2692 37092 2694
rect 37116 2692 37172 2694
rect 37196 2692 37252 2694
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 7616 2202 7672 2204
rect 7696 2202 7752 2204
rect 7776 2202 7832 2204
rect 7856 2202 7912 2204
rect 7616 2150 7662 2202
rect 7662 2150 7672 2202
rect 7696 2150 7726 2202
rect 7726 2150 7738 2202
rect 7738 2150 7752 2202
rect 7776 2150 7790 2202
rect 7790 2150 7802 2202
rect 7802 2150 7832 2202
rect 7856 2150 7866 2202
rect 7866 2150 7912 2202
rect 7616 2148 7672 2150
rect 7696 2148 7752 2150
rect 7776 2148 7832 2150
rect 7856 2148 7912 2150
rect 12616 2202 12672 2204
rect 12696 2202 12752 2204
rect 12776 2202 12832 2204
rect 12856 2202 12912 2204
rect 12616 2150 12662 2202
rect 12662 2150 12672 2202
rect 12696 2150 12726 2202
rect 12726 2150 12738 2202
rect 12738 2150 12752 2202
rect 12776 2150 12790 2202
rect 12790 2150 12802 2202
rect 12802 2150 12832 2202
rect 12856 2150 12866 2202
rect 12866 2150 12912 2202
rect 12616 2148 12672 2150
rect 12696 2148 12752 2150
rect 12776 2148 12832 2150
rect 12856 2148 12912 2150
rect 17616 2202 17672 2204
rect 17696 2202 17752 2204
rect 17776 2202 17832 2204
rect 17856 2202 17912 2204
rect 17616 2150 17662 2202
rect 17662 2150 17672 2202
rect 17696 2150 17726 2202
rect 17726 2150 17738 2202
rect 17738 2150 17752 2202
rect 17776 2150 17790 2202
rect 17790 2150 17802 2202
rect 17802 2150 17832 2202
rect 17856 2150 17866 2202
rect 17866 2150 17912 2202
rect 17616 2148 17672 2150
rect 17696 2148 17752 2150
rect 17776 2148 17832 2150
rect 17856 2148 17912 2150
rect 22616 2202 22672 2204
rect 22696 2202 22752 2204
rect 22776 2202 22832 2204
rect 22856 2202 22912 2204
rect 22616 2150 22662 2202
rect 22662 2150 22672 2202
rect 22696 2150 22726 2202
rect 22726 2150 22738 2202
rect 22738 2150 22752 2202
rect 22776 2150 22790 2202
rect 22790 2150 22802 2202
rect 22802 2150 22832 2202
rect 22856 2150 22866 2202
rect 22866 2150 22912 2202
rect 22616 2148 22672 2150
rect 22696 2148 22752 2150
rect 22776 2148 22832 2150
rect 22856 2148 22912 2150
rect 27616 2202 27672 2204
rect 27696 2202 27752 2204
rect 27776 2202 27832 2204
rect 27856 2202 27912 2204
rect 27616 2150 27662 2202
rect 27662 2150 27672 2202
rect 27696 2150 27726 2202
rect 27726 2150 27738 2202
rect 27738 2150 27752 2202
rect 27776 2150 27790 2202
rect 27790 2150 27802 2202
rect 27802 2150 27832 2202
rect 27856 2150 27866 2202
rect 27866 2150 27912 2202
rect 27616 2148 27672 2150
rect 27696 2148 27752 2150
rect 27776 2148 27832 2150
rect 27856 2148 27912 2150
rect 32616 2202 32672 2204
rect 32696 2202 32752 2204
rect 32776 2202 32832 2204
rect 32856 2202 32912 2204
rect 32616 2150 32662 2202
rect 32662 2150 32672 2202
rect 32696 2150 32726 2202
rect 32726 2150 32738 2202
rect 32738 2150 32752 2202
rect 32776 2150 32790 2202
rect 32790 2150 32802 2202
rect 32802 2150 32832 2202
rect 32856 2150 32866 2202
rect 32866 2150 32912 2202
rect 32616 2148 32672 2150
rect 32696 2148 32752 2150
rect 32776 2148 32832 2150
rect 32856 2148 32912 2150
rect 37616 2202 37672 2204
rect 37696 2202 37752 2204
rect 37776 2202 37832 2204
rect 37856 2202 37912 2204
rect 37616 2150 37662 2202
rect 37662 2150 37672 2202
rect 37696 2150 37726 2202
rect 37726 2150 37738 2202
rect 37738 2150 37752 2202
rect 37776 2150 37790 2202
rect 37790 2150 37802 2202
rect 37802 2150 37832 2202
rect 37856 2150 37866 2202
rect 37866 2150 37912 2202
rect 37616 2148 37672 2150
rect 37696 2148 37752 2150
rect 37776 2148 37832 2150
rect 37856 2148 37912 2150
<< metal3 >>
rect 1946 37568 2262 37569
rect 1946 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2262 37568
rect 1946 37503 2262 37504
rect 6946 37568 7262 37569
rect 6946 37504 6952 37568
rect 7016 37504 7032 37568
rect 7096 37504 7112 37568
rect 7176 37504 7192 37568
rect 7256 37504 7262 37568
rect 6946 37503 7262 37504
rect 11946 37568 12262 37569
rect 11946 37504 11952 37568
rect 12016 37504 12032 37568
rect 12096 37504 12112 37568
rect 12176 37504 12192 37568
rect 12256 37504 12262 37568
rect 11946 37503 12262 37504
rect 16946 37568 17262 37569
rect 16946 37504 16952 37568
rect 17016 37504 17032 37568
rect 17096 37504 17112 37568
rect 17176 37504 17192 37568
rect 17256 37504 17262 37568
rect 16946 37503 17262 37504
rect 21946 37568 22262 37569
rect 21946 37504 21952 37568
rect 22016 37504 22032 37568
rect 22096 37504 22112 37568
rect 22176 37504 22192 37568
rect 22256 37504 22262 37568
rect 21946 37503 22262 37504
rect 26946 37568 27262 37569
rect 26946 37504 26952 37568
rect 27016 37504 27032 37568
rect 27096 37504 27112 37568
rect 27176 37504 27192 37568
rect 27256 37504 27262 37568
rect 26946 37503 27262 37504
rect 31946 37568 32262 37569
rect 31946 37504 31952 37568
rect 32016 37504 32032 37568
rect 32096 37504 32112 37568
rect 32176 37504 32192 37568
rect 32256 37504 32262 37568
rect 31946 37503 32262 37504
rect 36946 37568 37262 37569
rect 36946 37504 36952 37568
rect 37016 37504 37032 37568
rect 37096 37504 37112 37568
rect 37176 37504 37192 37568
rect 37256 37504 37262 37568
rect 36946 37503 37262 37504
rect 2606 37024 2922 37025
rect 2606 36960 2612 37024
rect 2676 36960 2692 37024
rect 2756 36960 2772 37024
rect 2836 36960 2852 37024
rect 2916 36960 2922 37024
rect 2606 36959 2922 36960
rect 7606 37024 7922 37025
rect 7606 36960 7612 37024
rect 7676 36960 7692 37024
rect 7756 36960 7772 37024
rect 7836 36960 7852 37024
rect 7916 36960 7922 37024
rect 7606 36959 7922 36960
rect 12606 37024 12922 37025
rect 12606 36960 12612 37024
rect 12676 36960 12692 37024
rect 12756 36960 12772 37024
rect 12836 36960 12852 37024
rect 12916 36960 12922 37024
rect 12606 36959 12922 36960
rect 17606 37024 17922 37025
rect 17606 36960 17612 37024
rect 17676 36960 17692 37024
rect 17756 36960 17772 37024
rect 17836 36960 17852 37024
rect 17916 36960 17922 37024
rect 17606 36959 17922 36960
rect 22606 37024 22922 37025
rect 22606 36960 22612 37024
rect 22676 36960 22692 37024
rect 22756 36960 22772 37024
rect 22836 36960 22852 37024
rect 22916 36960 22922 37024
rect 22606 36959 22922 36960
rect 27606 37024 27922 37025
rect 27606 36960 27612 37024
rect 27676 36960 27692 37024
rect 27756 36960 27772 37024
rect 27836 36960 27852 37024
rect 27916 36960 27922 37024
rect 27606 36959 27922 36960
rect 32606 37024 32922 37025
rect 32606 36960 32612 37024
rect 32676 36960 32692 37024
rect 32756 36960 32772 37024
rect 32836 36960 32852 37024
rect 32916 36960 32922 37024
rect 32606 36959 32922 36960
rect 37606 37024 37922 37025
rect 37606 36960 37612 37024
rect 37676 36960 37692 37024
rect 37756 36960 37772 37024
rect 37836 36960 37852 37024
rect 37916 36960 37922 37024
rect 37606 36959 37922 36960
rect 1946 36480 2262 36481
rect 1946 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2262 36480
rect 1946 36415 2262 36416
rect 6946 36480 7262 36481
rect 6946 36416 6952 36480
rect 7016 36416 7032 36480
rect 7096 36416 7112 36480
rect 7176 36416 7192 36480
rect 7256 36416 7262 36480
rect 6946 36415 7262 36416
rect 11946 36480 12262 36481
rect 11946 36416 11952 36480
rect 12016 36416 12032 36480
rect 12096 36416 12112 36480
rect 12176 36416 12192 36480
rect 12256 36416 12262 36480
rect 11946 36415 12262 36416
rect 16946 36480 17262 36481
rect 16946 36416 16952 36480
rect 17016 36416 17032 36480
rect 17096 36416 17112 36480
rect 17176 36416 17192 36480
rect 17256 36416 17262 36480
rect 16946 36415 17262 36416
rect 21946 36480 22262 36481
rect 21946 36416 21952 36480
rect 22016 36416 22032 36480
rect 22096 36416 22112 36480
rect 22176 36416 22192 36480
rect 22256 36416 22262 36480
rect 21946 36415 22262 36416
rect 26946 36480 27262 36481
rect 26946 36416 26952 36480
rect 27016 36416 27032 36480
rect 27096 36416 27112 36480
rect 27176 36416 27192 36480
rect 27256 36416 27262 36480
rect 26946 36415 27262 36416
rect 31946 36480 32262 36481
rect 31946 36416 31952 36480
rect 32016 36416 32032 36480
rect 32096 36416 32112 36480
rect 32176 36416 32192 36480
rect 32256 36416 32262 36480
rect 31946 36415 32262 36416
rect 36946 36480 37262 36481
rect 36946 36416 36952 36480
rect 37016 36416 37032 36480
rect 37096 36416 37112 36480
rect 37176 36416 37192 36480
rect 37256 36416 37262 36480
rect 36946 36415 37262 36416
rect 2606 35936 2922 35937
rect 2606 35872 2612 35936
rect 2676 35872 2692 35936
rect 2756 35872 2772 35936
rect 2836 35872 2852 35936
rect 2916 35872 2922 35936
rect 2606 35871 2922 35872
rect 7606 35936 7922 35937
rect 7606 35872 7612 35936
rect 7676 35872 7692 35936
rect 7756 35872 7772 35936
rect 7836 35872 7852 35936
rect 7916 35872 7922 35936
rect 7606 35871 7922 35872
rect 12606 35936 12922 35937
rect 12606 35872 12612 35936
rect 12676 35872 12692 35936
rect 12756 35872 12772 35936
rect 12836 35872 12852 35936
rect 12916 35872 12922 35936
rect 12606 35871 12922 35872
rect 17606 35936 17922 35937
rect 17606 35872 17612 35936
rect 17676 35872 17692 35936
rect 17756 35872 17772 35936
rect 17836 35872 17852 35936
rect 17916 35872 17922 35936
rect 17606 35871 17922 35872
rect 22606 35936 22922 35937
rect 22606 35872 22612 35936
rect 22676 35872 22692 35936
rect 22756 35872 22772 35936
rect 22836 35872 22852 35936
rect 22916 35872 22922 35936
rect 22606 35871 22922 35872
rect 27606 35936 27922 35937
rect 27606 35872 27612 35936
rect 27676 35872 27692 35936
rect 27756 35872 27772 35936
rect 27836 35872 27852 35936
rect 27916 35872 27922 35936
rect 27606 35871 27922 35872
rect 32606 35936 32922 35937
rect 32606 35872 32612 35936
rect 32676 35872 32692 35936
rect 32756 35872 32772 35936
rect 32836 35872 32852 35936
rect 32916 35872 32922 35936
rect 32606 35871 32922 35872
rect 37606 35936 37922 35937
rect 37606 35872 37612 35936
rect 37676 35872 37692 35936
rect 37756 35872 37772 35936
rect 37836 35872 37852 35936
rect 37916 35872 37922 35936
rect 37606 35871 37922 35872
rect 1946 35392 2262 35393
rect 1946 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2262 35392
rect 1946 35327 2262 35328
rect 6946 35392 7262 35393
rect 6946 35328 6952 35392
rect 7016 35328 7032 35392
rect 7096 35328 7112 35392
rect 7176 35328 7192 35392
rect 7256 35328 7262 35392
rect 6946 35327 7262 35328
rect 11946 35392 12262 35393
rect 11946 35328 11952 35392
rect 12016 35328 12032 35392
rect 12096 35328 12112 35392
rect 12176 35328 12192 35392
rect 12256 35328 12262 35392
rect 11946 35327 12262 35328
rect 16946 35392 17262 35393
rect 16946 35328 16952 35392
rect 17016 35328 17032 35392
rect 17096 35328 17112 35392
rect 17176 35328 17192 35392
rect 17256 35328 17262 35392
rect 16946 35327 17262 35328
rect 21946 35392 22262 35393
rect 21946 35328 21952 35392
rect 22016 35328 22032 35392
rect 22096 35328 22112 35392
rect 22176 35328 22192 35392
rect 22256 35328 22262 35392
rect 21946 35327 22262 35328
rect 26946 35392 27262 35393
rect 26946 35328 26952 35392
rect 27016 35328 27032 35392
rect 27096 35328 27112 35392
rect 27176 35328 27192 35392
rect 27256 35328 27262 35392
rect 26946 35327 27262 35328
rect 31946 35392 32262 35393
rect 31946 35328 31952 35392
rect 32016 35328 32032 35392
rect 32096 35328 32112 35392
rect 32176 35328 32192 35392
rect 32256 35328 32262 35392
rect 31946 35327 32262 35328
rect 36946 35392 37262 35393
rect 36946 35328 36952 35392
rect 37016 35328 37032 35392
rect 37096 35328 37112 35392
rect 37176 35328 37192 35392
rect 37256 35328 37262 35392
rect 36946 35327 37262 35328
rect 2606 34848 2922 34849
rect 2606 34784 2612 34848
rect 2676 34784 2692 34848
rect 2756 34784 2772 34848
rect 2836 34784 2852 34848
rect 2916 34784 2922 34848
rect 2606 34783 2922 34784
rect 7606 34848 7922 34849
rect 7606 34784 7612 34848
rect 7676 34784 7692 34848
rect 7756 34784 7772 34848
rect 7836 34784 7852 34848
rect 7916 34784 7922 34848
rect 7606 34783 7922 34784
rect 12606 34848 12922 34849
rect 12606 34784 12612 34848
rect 12676 34784 12692 34848
rect 12756 34784 12772 34848
rect 12836 34784 12852 34848
rect 12916 34784 12922 34848
rect 12606 34783 12922 34784
rect 17606 34848 17922 34849
rect 17606 34784 17612 34848
rect 17676 34784 17692 34848
rect 17756 34784 17772 34848
rect 17836 34784 17852 34848
rect 17916 34784 17922 34848
rect 17606 34783 17922 34784
rect 22606 34848 22922 34849
rect 22606 34784 22612 34848
rect 22676 34784 22692 34848
rect 22756 34784 22772 34848
rect 22836 34784 22852 34848
rect 22916 34784 22922 34848
rect 22606 34783 22922 34784
rect 27606 34848 27922 34849
rect 27606 34784 27612 34848
rect 27676 34784 27692 34848
rect 27756 34784 27772 34848
rect 27836 34784 27852 34848
rect 27916 34784 27922 34848
rect 27606 34783 27922 34784
rect 32606 34848 32922 34849
rect 32606 34784 32612 34848
rect 32676 34784 32692 34848
rect 32756 34784 32772 34848
rect 32836 34784 32852 34848
rect 32916 34784 32922 34848
rect 32606 34783 32922 34784
rect 37606 34848 37922 34849
rect 37606 34784 37612 34848
rect 37676 34784 37692 34848
rect 37756 34784 37772 34848
rect 37836 34784 37852 34848
rect 37916 34784 37922 34848
rect 37606 34783 37922 34784
rect 1946 34304 2262 34305
rect 1946 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2262 34304
rect 1946 34239 2262 34240
rect 6946 34304 7262 34305
rect 6946 34240 6952 34304
rect 7016 34240 7032 34304
rect 7096 34240 7112 34304
rect 7176 34240 7192 34304
rect 7256 34240 7262 34304
rect 6946 34239 7262 34240
rect 11946 34304 12262 34305
rect 11946 34240 11952 34304
rect 12016 34240 12032 34304
rect 12096 34240 12112 34304
rect 12176 34240 12192 34304
rect 12256 34240 12262 34304
rect 11946 34239 12262 34240
rect 16946 34304 17262 34305
rect 16946 34240 16952 34304
rect 17016 34240 17032 34304
rect 17096 34240 17112 34304
rect 17176 34240 17192 34304
rect 17256 34240 17262 34304
rect 16946 34239 17262 34240
rect 21946 34304 22262 34305
rect 21946 34240 21952 34304
rect 22016 34240 22032 34304
rect 22096 34240 22112 34304
rect 22176 34240 22192 34304
rect 22256 34240 22262 34304
rect 21946 34239 22262 34240
rect 26946 34304 27262 34305
rect 26946 34240 26952 34304
rect 27016 34240 27032 34304
rect 27096 34240 27112 34304
rect 27176 34240 27192 34304
rect 27256 34240 27262 34304
rect 26946 34239 27262 34240
rect 31946 34304 32262 34305
rect 31946 34240 31952 34304
rect 32016 34240 32032 34304
rect 32096 34240 32112 34304
rect 32176 34240 32192 34304
rect 32256 34240 32262 34304
rect 31946 34239 32262 34240
rect 36946 34304 37262 34305
rect 36946 34240 36952 34304
rect 37016 34240 37032 34304
rect 37096 34240 37112 34304
rect 37176 34240 37192 34304
rect 37256 34240 37262 34304
rect 36946 34239 37262 34240
rect 2606 33760 2922 33761
rect 2606 33696 2612 33760
rect 2676 33696 2692 33760
rect 2756 33696 2772 33760
rect 2836 33696 2852 33760
rect 2916 33696 2922 33760
rect 2606 33695 2922 33696
rect 7606 33760 7922 33761
rect 7606 33696 7612 33760
rect 7676 33696 7692 33760
rect 7756 33696 7772 33760
rect 7836 33696 7852 33760
rect 7916 33696 7922 33760
rect 7606 33695 7922 33696
rect 12606 33760 12922 33761
rect 12606 33696 12612 33760
rect 12676 33696 12692 33760
rect 12756 33696 12772 33760
rect 12836 33696 12852 33760
rect 12916 33696 12922 33760
rect 12606 33695 12922 33696
rect 17606 33760 17922 33761
rect 17606 33696 17612 33760
rect 17676 33696 17692 33760
rect 17756 33696 17772 33760
rect 17836 33696 17852 33760
rect 17916 33696 17922 33760
rect 17606 33695 17922 33696
rect 22606 33760 22922 33761
rect 22606 33696 22612 33760
rect 22676 33696 22692 33760
rect 22756 33696 22772 33760
rect 22836 33696 22852 33760
rect 22916 33696 22922 33760
rect 22606 33695 22922 33696
rect 27606 33760 27922 33761
rect 27606 33696 27612 33760
rect 27676 33696 27692 33760
rect 27756 33696 27772 33760
rect 27836 33696 27852 33760
rect 27916 33696 27922 33760
rect 27606 33695 27922 33696
rect 32606 33760 32922 33761
rect 32606 33696 32612 33760
rect 32676 33696 32692 33760
rect 32756 33696 32772 33760
rect 32836 33696 32852 33760
rect 32916 33696 32922 33760
rect 32606 33695 32922 33696
rect 37606 33760 37922 33761
rect 37606 33696 37612 33760
rect 37676 33696 37692 33760
rect 37756 33696 37772 33760
rect 37836 33696 37852 33760
rect 37916 33696 37922 33760
rect 37606 33695 37922 33696
rect 1946 33216 2262 33217
rect 1946 33152 1952 33216
rect 2016 33152 2032 33216
rect 2096 33152 2112 33216
rect 2176 33152 2192 33216
rect 2256 33152 2262 33216
rect 1946 33151 2262 33152
rect 6946 33216 7262 33217
rect 6946 33152 6952 33216
rect 7016 33152 7032 33216
rect 7096 33152 7112 33216
rect 7176 33152 7192 33216
rect 7256 33152 7262 33216
rect 6946 33151 7262 33152
rect 11946 33216 12262 33217
rect 11946 33152 11952 33216
rect 12016 33152 12032 33216
rect 12096 33152 12112 33216
rect 12176 33152 12192 33216
rect 12256 33152 12262 33216
rect 11946 33151 12262 33152
rect 16946 33216 17262 33217
rect 16946 33152 16952 33216
rect 17016 33152 17032 33216
rect 17096 33152 17112 33216
rect 17176 33152 17192 33216
rect 17256 33152 17262 33216
rect 16946 33151 17262 33152
rect 21946 33216 22262 33217
rect 21946 33152 21952 33216
rect 22016 33152 22032 33216
rect 22096 33152 22112 33216
rect 22176 33152 22192 33216
rect 22256 33152 22262 33216
rect 21946 33151 22262 33152
rect 26946 33216 27262 33217
rect 26946 33152 26952 33216
rect 27016 33152 27032 33216
rect 27096 33152 27112 33216
rect 27176 33152 27192 33216
rect 27256 33152 27262 33216
rect 26946 33151 27262 33152
rect 31946 33216 32262 33217
rect 31946 33152 31952 33216
rect 32016 33152 32032 33216
rect 32096 33152 32112 33216
rect 32176 33152 32192 33216
rect 32256 33152 32262 33216
rect 31946 33151 32262 33152
rect 36946 33216 37262 33217
rect 36946 33152 36952 33216
rect 37016 33152 37032 33216
rect 37096 33152 37112 33216
rect 37176 33152 37192 33216
rect 37256 33152 37262 33216
rect 36946 33151 37262 33152
rect 2606 32672 2922 32673
rect 2606 32608 2612 32672
rect 2676 32608 2692 32672
rect 2756 32608 2772 32672
rect 2836 32608 2852 32672
rect 2916 32608 2922 32672
rect 2606 32607 2922 32608
rect 7606 32672 7922 32673
rect 7606 32608 7612 32672
rect 7676 32608 7692 32672
rect 7756 32608 7772 32672
rect 7836 32608 7852 32672
rect 7916 32608 7922 32672
rect 7606 32607 7922 32608
rect 12606 32672 12922 32673
rect 12606 32608 12612 32672
rect 12676 32608 12692 32672
rect 12756 32608 12772 32672
rect 12836 32608 12852 32672
rect 12916 32608 12922 32672
rect 12606 32607 12922 32608
rect 17606 32672 17922 32673
rect 17606 32608 17612 32672
rect 17676 32608 17692 32672
rect 17756 32608 17772 32672
rect 17836 32608 17852 32672
rect 17916 32608 17922 32672
rect 17606 32607 17922 32608
rect 22606 32672 22922 32673
rect 22606 32608 22612 32672
rect 22676 32608 22692 32672
rect 22756 32608 22772 32672
rect 22836 32608 22852 32672
rect 22916 32608 22922 32672
rect 22606 32607 22922 32608
rect 27606 32672 27922 32673
rect 27606 32608 27612 32672
rect 27676 32608 27692 32672
rect 27756 32608 27772 32672
rect 27836 32608 27852 32672
rect 27916 32608 27922 32672
rect 27606 32607 27922 32608
rect 32606 32672 32922 32673
rect 32606 32608 32612 32672
rect 32676 32608 32692 32672
rect 32756 32608 32772 32672
rect 32836 32608 32852 32672
rect 32916 32608 32922 32672
rect 32606 32607 32922 32608
rect 37606 32672 37922 32673
rect 37606 32608 37612 32672
rect 37676 32608 37692 32672
rect 37756 32608 37772 32672
rect 37836 32608 37852 32672
rect 37916 32608 37922 32672
rect 37606 32607 37922 32608
rect 1946 32128 2262 32129
rect 1946 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2262 32128
rect 1946 32063 2262 32064
rect 6946 32128 7262 32129
rect 6946 32064 6952 32128
rect 7016 32064 7032 32128
rect 7096 32064 7112 32128
rect 7176 32064 7192 32128
rect 7256 32064 7262 32128
rect 6946 32063 7262 32064
rect 11946 32128 12262 32129
rect 11946 32064 11952 32128
rect 12016 32064 12032 32128
rect 12096 32064 12112 32128
rect 12176 32064 12192 32128
rect 12256 32064 12262 32128
rect 11946 32063 12262 32064
rect 16946 32128 17262 32129
rect 16946 32064 16952 32128
rect 17016 32064 17032 32128
rect 17096 32064 17112 32128
rect 17176 32064 17192 32128
rect 17256 32064 17262 32128
rect 16946 32063 17262 32064
rect 21946 32128 22262 32129
rect 21946 32064 21952 32128
rect 22016 32064 22032 32128
rect 22096 32064 22112 32128
rect 22176 32064 22192 32128
rect 22256 32064 22262 32128
rect 21946 32063 22262 32064
rect 26946 32128 27262 32129
rect 26946 32064 26952 32128
rect 27016 32064 27032 32128
rect 27096 32064 27112 32128
rect 27176 32064 27192 32128
rect 27256 32064 27262 32128
rect 26946 32063 27262 32064
rect 31946 32128 32262 32129
rect 31946 32064 31952 32128
rect 32016 32064 32032 32128
rect 32096 32064 32112 32128
rect 32176 32064 32192 32128
rect 32256 32064 32262 32128
rect 31946 32063 32262 32064
rect 36946 32128 37262 32129
rect 36946 32064 36952 32128
rect 37016 32064 37032 32128
rect 37096 32064 37112 32128
rect 37176 32064 37192 32128
rect 37256 32064 37262 32128
rect 36946 32063 37262 32064
rect 2606 31584 2922 31585
rect 2606 31520 2612 31584
rect 2676 31520 2692 31584
rect 2756 31520 2772 31584
rect 2836 31520 2852 31584
rect 2916 31520 2922 31584
rect 2606 31519 2922 31520
rect 7606 31584 7922 31585
rect 7606 31520 7612 31584
rect 7676 31520 7692 31584
rect 7756 31520 7772 31584
rect 7836 31520 7852 31584
rect 7916 31520 7922 31584
rect 7606 31519 7922 31520
rect 12606 31584 12922 31585
rect 12606 31520 12612 31584
rect 12676 31520 12692 31584
rect 12756 31520 12772 31584
rect 12836 31520 12852 31584
rect 12916 31520 12922 31584
rect 12606 31519 12922 31520
rect 17606 31584 17922 31585
rect 17606 31520 17612 31584
rect 17676 31520 17692 31584
rect 17756 31520 17772 31584
rect 17836 31520 17852 31584
rect 17916 31520 17922 31584
rect 17606 31519 17922 31520
rect 22606 31584 22922 31585
rect 22606 31520 22612 31584
rect 22676 31520 22692 31584
rect 22756 31520 22772 31584
rect 22836 31520 22852 31584
rect 22916 31520 22922 31584
rect 22606 31519 22922 31520
rect 27606 31584 27922 31585
rect 27606 31520 27612 31584
rect 27676 31520 27692 31584
rect 27756 31520 27772 31584
rect 27836 31520 27852 31584
rect 27916 31520 27922 31584
rect 27606 31519 27922 31520
rect 32606 31584 32922 31585
rect 32606 31520 32612 31584
rect 32676 31520 32692 31584
rect 32756 31520 32772 31584
rect 32836 31520 32852 31584
rect 32916 31520 32922 31584
rect 32606 31519 32922 31520
rect 37606 31584 37922 31585
rect 37606 31520 37612 31584
rect 37676 31520 37692 31584
rect 37756 31520 37772 31584
rect 37836 31520 37852 31584
rect 37916 31520 37922 31584
rect 37606 31519 37922 31520
rect 1946 31040 2262 31041
rect 1946 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2262 31040
rect 1946 30975 2262 30976
rect 6946 31040 7262 31041
rect 6946 30976 6952 31040
rect 7016 30976 7032 31040
rect 7096 30976 7112 31040
rect 7176 30976 7192 31040
rect 7256 30976 7262 31040
rect 6946 30975 7262 30976
rect 11946 31040 12262 31041
rect 11946 30976 11952 31040
rect 12016 30976 12032 31040
rect 12096 30976 12112 31040
rect 12176 30976 12192 31040
rect 12256 30976 12262 31040
rect 11946 30975 12262 30976
rect 16946 31040 17262 31041
rect 16946 30976 16952 31040
rect 17016 30976 17032 31040
rect 17096 30976 17112 31040
rect 17176 30976 17192 31040
rect 17256 30976 17262 31040
rect 16946 30975 17262 30976
rect 21946 31040 22262 31041
rect 21946 30976 21952 31040
rect 22016 30976 22032 31040
rect 22096 30976 22112 31040
rect 22176 30976 22192 31040
rect 22256 30976 22262 31040
rect 21946 30975 22262 30976
rect 26946 31040 27262 31041
rect 26946 30976 26952 31040
rect 27016 30976 27032 31040
rect 27096 30976 27112 31040
rect 27176 30976 27192 31040
rect 27256 30976 27262 31040
rect 26946 30975 27262 30976
rect 31946 31040 32262 31041
rect 31946 30976 31952 31040
rect 32016 30976 32032 31040
rect 32096 30976 32112 31040
rect 32176 30976 32192 31040
rect 32256 30976 32262 31040
rect 31946 30975 32262 30976
rect 36946 31040 37262 31041
rect 36946 30976 36952 31040
rect 37016 30976 37032 31040
rect 37096 30976 37112 31040
rect 37176 30976 37192 31040
rect 37256 30976 37262 31040
rect 36946 30975 37262 30976
rect 2606 30496 2922 30497
rect 2606 30432 2612 30496
rect 2676 30432 2692 30496
rect 2756 30432 2772 30496
rect 2836 30432 2852 30496
rect 2916 30432 2922 30496
rect 2606 30431 2922 30432
rect 7606 30496 7922 30497
rect 7606 30432 7612 30496
rect 7676 30432 7692 30496
rect 7756 30432 7772 30496
rect 7836 30432 7852 30496
rect 7916 30432 7922 30496
rect 7606 30431 7922 30432
rect 12606 30496 12922 30497
rect 12606 30432 12612 30496
rect 12676 30432 12692 30496
rect 12756 30432 12772 30496
rect 12836 30432 12852 30496
rect 12916 30432 12922 30496
rect 12606 30431 12922 30432
rect 17606 30496 17922 30497
rect 17606 30432 17612 30496
rect 17676 30432 17692 30496
rect 17756 30432 17772 30496
rect 17836 30432 17852 30496
rect 17916 30432 17922 30496
rect 17606 30431 17922 30432
rect 22606 30496 22922 30497
rect 22606 30432 22612 30496
rect 22676 30432 22692 30496
rect 22756 30432 22772 30496
rect 22836 30432 22852 30496
rect 22916 30432 22922 30496
rect 22606 30431 22922 30432
rect 27606 30496 27922 30497
rect 27606 30432 27612 30496
rect 27676 30432 27692 30496
rect 27756 30432 27772 30496
rect 27836 30432 27852 30496
rect 27916 30432 27922 30496
rect 27606 30431 27922 30432
rect 32606 30496 32922 30497
rect 32606 30432 32612 30496
rect 32676 30432 32692 30496
rect 32756 30432 32772 30496
rect 32836 30432 32852 30496
rect 32916 30432 32922 30496
rect 32606 30431 32922 30432
rect 37606 30496 37922 30497
rect 37606 30432 37612 30496
rect 37676 30432 37692 30496
rect 37756 30432 37772 30496
rect 37836 30432 37852 30496
rect 37916 30432 37922 30496
rect 37606 30431 37922 30432
rect 1946 29952 2262 29953
rect 1946 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2262 29952
rect 1946 29887 2262 29888
rect 6946 29952 7262 29953
rect 6946 29888 6952 29952
rect 7016 29888 7032 29952
rect 7096 29888 7112 29952
rect 7176 29888 7192 29952
rect 7256 29888 7262 29952
rect 6946 29887 7262 29888
rect 11946 29952 12262 29953
rect 11946 29888 11952 29952
rect 12016 29888 12032 29952
rect 12096 29888 12112 29952
rect 12176 29888 12192 29952
rect 12256 29888 12262 29952
rect 11946 29887 12262 29888
rect 16946 29952 17262 29953
rect 16946 29888 16952 29952
rect 17016 29888 17032 29952
rect 17096 29888 17112 29952
rect 17176 29888 17192 29952
rect 17256 29888 17262 29952
rect 16946 29887 17262 29888
rect 21946 29952 22262 29953
rect 21946 29888 21952 29952
rect 22016 29888 22032 29952
rect 22096 29888 22112 29952
rect 22176 29888 22192 29952
rect 22256 29888 22262 29952
rect 21946 29887 22262 29888
rect 26946 29952 27262 29953
rect 26946 29888 26952 29952
rect 27016 29888 27032 29952
rect 27096 29888 27112 29952
rect 27176 29888 27192 29952
rect 27256 29888 27262 29952
rect 26946 29887 27262 29888
rect 31946 29952 32262 29953
rect 31946 29888 31952 29952
rect 32016 29888 32032 29952
rect 32096 29888 32112 29952
rect 32176 29888 32192 29952
rect 32256 29888 32262 29952
rect 31946 29887 32262 29888
rect 36946 29952 37262 29953
rect 36946 29888 36952 29952
rect 37016 29888 37032 29952
rect 37096 29888 37112 29952
rect 37176 29888 37192 29952
rect 37256 29888 37262 29952
rect 36946 29887 37262 29888
rect 2606 29408 2922 29409
rect 2606 29344 2612 29408
rect 2676 29344 2692 29408
rect 2756 29344 2772 29408
rect 2836 29344 2852 29408
rect 2916 29344 2922 29408
rect 2606 29343 2922 29344
rect 7606 29408 7922 29409
rect 7606 29344 7612 29408
rect 7676 29344 7692 29408
rect 7756 29344 7772 29408
rect 7836 29344 7852 29408
rect 7916 29344 7922 29408
rect 7606 29343 7922 29344
rect 12606 29408 12922 29409
rect 12606 29344 12612 29408
rect 12676 29344 12692 29408
rect 12756 29344 12772 29408
rect 12836 29344 12852 29408
rect 12916 29344 12922 29408
rect 12606 29343 12922 29344
rect 17606 29408 17922 29409
rect 17606 29344 17612 29408
rect 17676 29344 17692 29408
rect 17756 29344 17772 29408
rect 17836 29344 17852 29408
rect 17916 29344 17922 29408
rect 17606 29343 17922 29344
rect 22606 29408 22922 29409
rect 22606 29344 22612 29408
rect 22676 29344 22692 29408
rect 22756 29344 22772 29408
rect 22836 29344 22852 29408
rect 22916 29344 22922 29408
rect 22606 29343 22922 29344
rect 27606 29408 27922 29409
rect 27606 29344 27612 29408
rect 27676 29344 27692 29408
rect 27756 29344 27772 29408
rect 27836 29344 27852 29408
rect 27916 29344 27922 29408
rect 27606 29343 27922 29344
rect 32606 29408 32922 29409
rect 32606 29344 32612 29408
rect 32676 29344 32692 29408
rect 32756 29344 32772 29408
rect 32836 29344 32852 29408
rect 32916 29344 32922 29408
rect 32606 29343 32922 29344
rect 37606 29408 37922 29409
rect 37606 29344 37612 29408
rect 37676 29344 37692 29408
rect 37756 29344 37772 29408
rect 37836 29344 37852 29408
rect 37916 29344 37922 29408
rect 37606 29343 37922 29344
rect 1946 28864 2262 28865
rect 1946 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2262 28864
rect 1946 28799 2262 28800
rect 6946 28864 7262 28865
rect 6946 28800 6952 28864
rect 7016 28800 7032 28864
rect 7096 28800 7112 28864
rect 7176 28800 7192 28864
rect 7256 28800 7262 28864
rect 6946 28799 7262 28800
rect 11946 28864 12262 28865
rect 11946 28800 11952 28864
rect 12016 28800 12032 28864
rect 12096 28800 12112 28864
rect 12176 28800 12192 28864
rect 12256 28800 12262 28864
rect 11946 28799 12262 28800
rect 16946 28864 17262 28865
rect 16946 28800 16952 28864
rect 17016 28800 17032 28864
rect 17096 28800 17112 28864
rect 17176 28800 17192 28864
rect 17256 28800 17262 28864
rect 16946 28799 17262 28800
rect 21946 28864 22262 28865
rect 21946 28800 21952 28864
rect 22016 28800 22032 28864
rect 22096 28800 22112 28864
rect 22176 28800 22192 28864
rect 22256 28800 22262 28864
rect 21946 28799 22262 28800
rect 26946 28864 27262 28865
rect 26946 28800 26952 28864
rect 27016 28800 27032 28864
rect 27096 28800 27112 28864
rect 27176 28800 27192 28864
rect 27256 28800 27262 28864
rect 26946 28799 27262 28800
rect 31946 28864 32262 28865
rect 31946 28800 31952 28864
rect 32016 28800 32032 28864
rect 32096 28800 32112 28864
rect 32176 28800 32192 28864
rect 32256 28800 32262 28864
rect 31946 28799 32262 28800
rect 36946 28864 37262 28865
rect 36946 28800 36952 28864
rect 37016 28800 37032 28864
rect 37096 28800 37112 28864
rect 37176 28800 37192 28864
rect 37256 28800 37262 28864
rect 36946 28799 37262 28800
rect 2606 28320 2922 28321
rect 2606 28256 2612 28320
rect 2676 28256 2692 28320
rect 2756 28256 2772 28320
rect 2836 28256 2852 28320
rect 2916 28256 2922 28320
rect 2606 28255 2922 28256
rect 7606 28320 7922 28321
rect 7606 28256 7612 28320
rect 7676 28256 7692 28320
rect 7756 28256 7772 28320
rect 7836 28256 7852 28320
rect 7916 28256 7922 28320
rect 7606 28255 7922 28256
rect 12606 28320 12922 28321
rect 12606 28256 12612 28320
rect 12676 28256 12692 28320
rect 12756 28256 12772 28320
rect 12836 28256 12852 28320
rect 12916 28256 12922 28320
rect 12606 28255 12922 28256
rect 17606 28320 17922 28321
rect 17606 28256 17612 28320
rect 17676 28256 17692 28320
rect 17756 28256 17772 28320
rect 17836 28256 17852 28320
rect 17916 28256 17922 28320
rect 17606 28255 17922 28256
rect 22606 28320 22922 28321
rect 22606 28256 22612 28320
rect 22676 28256 22692 28320
rect 22756 28256 22772 28320
rect 22836 28256 22852 28320
rect 22916 28256 22922 28320
rect 22606 28255 22922 28256
rect 27606 28320 27922 28321
rect 27606 28256 27612 28320
rect 27676 28256 27692 28320
rect 27756 28256 27772 28320
rect 27836 28256 27852 28320
rect 27916 28256 27922 28320
rect 27606 28255 27922 28256
rect 32606 28320 32922 28321
rect 32606 28256 32612 28320
rect 32676 28256 32692 28320
rect 32756 28256 32772 28320
rect 32836 28256 32852 28320
rect 32916 28256 32922 28320
rect 32606 28255 32922 28256
rect 37606 28320 37922 28321
rect 37606 28256 37612 28320
rect 37676 28256 37692 28320
rect 37756 28256 37772 28320
rect 37836 28256 37852 28320
rect 37916 28256 37922 28320
rect 37606 28255 37922 28256
rect 1946 27776 2262 27777
rect 1946 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2262 27776
rect 1946 27711 2262 27712
rect 6946 27776 7262 27777
rect 6946 27712 6952 27776
rect 7016 27712 7032 27776
rect 7096 27712 7112 27776
rect 7176 27712 7192 27776
rect 7256 27712 7262 27776
rect 6946 27711 7262 27712
rect 11946 27776 12262 27777
rect 11946 27712 11952 27776
rect 12016 27712 12032 27776
rect 12096 27712 12112 27776
rect 12176 27712 12192 27776
rect 12256 27712 12262 27776
rect 11946 27711 12262 27712
rect 16946 27776 17262 27777
rect 16946 27712 16952 27776
rect 17016 27712 17032 27776
rect 17096 27712 17112 27776
rect 17176 27712 17192 27776
rect 17256 27712 17262 27776
rect 16946 27711 17262 27712
rect 21946 27776 22262 27777
rect 21946 27712 21952 27776
rect 22016 27712 22032 27776
rect 22096 27712 22112 27776
rect 22176 27712 22192 27776
rect 22256 27712 22262 27776
rect 21946 27711 22262 27712
rect 26946 27776 27262 27777
rect 26946 27712 26952 27776
rect 27016 27712 27032 27776
rect 27096 27712 27112 27776
rect 27176 27712 27192 27776
rect 27256 27712 27262 27776
rect 26946 27711 27262 27712
rect 31946 27776 32262 27777
rect 31946 27712 31952 27776
rect 32016 27712 32032 27776
rect 32096 27712 32112 27776
rect 32176 27712 32192 27776
rect 32256 27712 32262 27776
rect 31946 27711 32262 27712
rect 36946 27776 37262 27777
rect 36946 27712 36952 27776
rect 37016 27712 37032 27776
rect 37096 27712 37112 27776
rect 37176 27712 37192 27776
rect 37256 27712 37262 27776
rect 36946 27711 37262 27712
rect 2606 27232 2922 27233
rect 2606 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2922 27232
rect 2606 27167 2922 27168
rect 7606 27232 7922 27233
rect 7606 27168 7612 27232
rect 7676 27168 7692 27232
rect 7756 27168 7772 27232
rect 7836 27168 7852 27232
rect 7916 27168 7922 27232
rect 7606 27167 7922 27168
rect 12606 27232 12922 27233
rect 12606 27168 12612 27232
rect 12676 27168 12692 27232
rect 12756 27168 12772 27232
rect 12836 27168 12852 27232
rect 12916 27168 12922 27232
rect 12606 27167 12922 27168
rect 17606 27232 17922 27233
rect 17606 27168 17612 27232
rect 17676 27168 17692 27232
rect 17756 27168 17772 27232
rect 17836 27168 17852 27232
rect 17916 27168 17922 27232
rect 17606 27167 17922 27168
rect 22606 27232 22922 27233
rect 22606 27168 22612 27232
rect 22676 27168 22692 27232
rect 22756 27168 22772 27232
rect 22836 27168 22852 27232
rect 22916 27168 22922 27232
rect 22606 27167 22922 27168
rect 27606 27232 27922 27233
rect 27606 27168 27612 27232
rect 27676 27168 27692 27232
rect 27756 27168 27772 27232
rect 27836 27168 27852 27232
rect 27916 27168 27922 27232
rect 27606 27167 27922 27168
rect 32606 27232 32922 27233
rect 32606 27168 32612 27232
rect 32676 27168 32692 27232
rect 32756 27168 32772 27232
rect 32836 27168 32852 27232
rect 32916 27168 32922 27232
rect 32606 27167 32922 27168
rect 37606 27232 37922 27233
rect 37606 27168 37612 27232
rect 37676 27168 37692 27232
rect 37756 27168 37772 27232
rect 37836 27168 37852 27232
rect 37916 27168 37922 27232
rect 37606 27167 37922 27168
rect 1946 26688 2262 26689
rect 1946 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2262 26688
rect 1946 26623 2262 26624
rect 6946 26688 7262 26689
rect 6946 26624 6952 26688
rect 7016 26624 7032 26688
rect 7096 26624 7112 26688
rect 7176 26624 7192 26688
rect 7256 26624 7262 26688
rect 6946 26623 7262 26624
rect 11946 26688 12262 26689
rect 11946 26624 11952 26688
rect 12016 26624 12032 26688
rect 12096 26624 12112 26688
rect 12176 26624 12192 26688
rect 12256 26624 12262 26688
rect 11946 26623 12262 26624
rect 16946 26688 17262 26689
rect 16946 26624 16952 26688
rect 17016 26624 17032 26688
rect 17096 26624 17112 26688
rect 17176 26624 17192 26688
rect 17256 26624 17262 26688
rect 16946 26623 17262 26624
rect 21946 26688 22262 26689
rect 21946 26624 21952 26688
rect 22016 26624 22032 26688
rect 22096 26624 22112 26688
rect 22176 26624 22192 26688
rect 22256 26624 22262 26688
rect 21946 26623 22262 26624
rect 26946 26688 27262 26689
rect 26946 26624 26952 26688
rect 27016 26624 27032 26688
rect 27096 26624 27112 26688
rect 27176 26624 27192 26688
rect 27256 26624 27262 26688
rect 26946 26623 27262 26624
rect 31946 26688 32262 26689
rect 31946 26624 31952 26688
rect 32016 26624 32032 26688
rect 32096 26624 32112 26688
rect 32176 26624 32192 26688
rect 32256 26624 32262 26688
rect 31946 26623 32262 26624
rect 36946 26688 37262 26689
rect 36946 26624 36952 26688
rect 37016 26624 37032 26688
rect 37096 26624 37112 26688
rect 37176 26624 37192 26688
rect 37256 26624 37262 26688
rect 36946 26623 37262 26624
rect 2606 26144 2922 26145
rect 2606 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2922 26144
rect 2606 26079 2922 26080
rect 7606 26144 7922 26145
rect 7606 26080 7612 26144
rect 7676 26080 7692 26144
rect 7756 26080 7772 26144
rect 7836 26080 7852 26144
rect 7916 26080 7922 26144
rect 7606 26079 7922 26080
rect 12606 26144 12922 26145
rect 12606 26080 12612 26144
rect 12676 26080 12692 26144
rect 12756 26080 12772 26144
rect 12836 26080 12852 26144
rect 12916 26080 12922 26144
rect 12606 26079 12922 26080
rect 17606 26144 17922 26145
rect 17606 26080 17612 26144
rect 17676 26080 17692 26144
rect 17756 26080 17772 26144
rect 17836 26080 17852 26144
rect 17916 26080 17922 26144
rect 17606 26079 17922 26080
rect 22606 26144 22922 26145
rect 22606 26080 22612 26144
rect 22676 26080 22692 26144
rect 22756 26080 22772 26144
rect 22836 26080 22852 26144
rect 22916 26080 22922 26144
rect 22606 26079 22922 26080
rect 27606 26144 27922 26145
rect 27606 26080 27612 26144
rect 27676 26080 27692 26144
rect 27756 26080 27772 26144
rect 27836 26080 27852 26144
rect 27916 26080 27922 26144
rect 27606 26079 27922 26080
rect 32606 26144 32922 26145
rect 32606 26080 32612 26144
rect 32676 26080 32692 26144
rect 32756 26080 32772 26144
rect 32836 26080 32852 26144
rect 32916 26080 32922 26144
rect 32606 26079 32922 26080
rect 37606 26144 37922 26145
rect 37606 26080 37612 26144
rect 37676 26080 37692 26144
rect 37756 26080 37772 26144
rect 37836 26080 37852 26144
rect 37916 26080 37922 26144
rect 37606 26079 37922 26080
rect 1946 25600 2262 25601
rect 1946 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2262 25600
rect 1946 25535 2262 25536
rect 6946 25600 7262 25601
rect 6946 25536 6952 25600
rect 7016 25536 7032 25600
rect 7096 25536 7112 25600
rect 7176 25536 7192 25600
rect 7256 25536 7262 25600
rect 6946 25535 7262 25536
rect 11946 25600 12262 25601
rect 11946 25536 11952 25600
rect 12016 25536 12032 25600
rect 12096 25536 12112 25600
rect 12176 25536 12192 25600
rect 12256 25536 12262 25600
rect 11946 25535 12262 25536
rect 16946 25600 17262 25601
rect 16946 25536 16952 25600
rect 17016 25536 17032 25600
rect 17096 25536 17112 25600
rect 17176 25536 17192 25600
rect 17256 25536 17262 25600
rect 16946 25535 17262 25536
rect 21946 25600 22262 25601
rect 21946 25536 21952 25600
rect 22016 25536 22032 25600
rect 22096 25536 22112 25600
rect 22176 25536 22192 25600
rect 22256 25536 22262 25600
rect 21946 25535 22262 25536
rect 26946 25600 27262 25601
rect 26946 25536 26952 25600
rect 27016 25536 27032 25600
rect 27096 25536 27112 25600
rect 27176 25536 27192 25600
rect 27256 25536 27262 25600
rect 26946 25535 27262 25536
rect 31946 25600 32262 25601
rect 31946 25536 31952 25600
rect 32016 25536 32032 25600
rect 32096 25536 32112 25600
rect 32176 25536 32192 25600
rect 32256 25536 32262 25600
rect 31946 25535 32262 25536
rect 36946 25600 37262 25601
rect 36946 25536 36952 25600
rect 37016 25536 37032 25600
rect 37096 25536 37112 25600
rect 37176 25536 37192 25600
rect 37256 25536 37262 25600
rect 36946 25535 37262 25536
rect 2606 25056 2922 25057
rect 2606 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2922 25056
rect 2606 24991 2922 24992
rect 7606 25056 7922 25057
rect 7606 24992 7612 25056
rect 7676 24992 7692 25056
rect 7756 24992 7772 25056
rect 7836 24992 7852 25056
rect 7916 24992 7922 25056
rect 7606 24991 7922 24992
rect 12606 25056 12922 25057
rect 12606 24992 12612 25056
rect 12676 24992 12692 25056
rect 12756 24992 12772 25056
rect 12836 24992 12852 25056
rect 12916 24992 12922 25056
rect 12606 24991 12922 24992
rect 17606 25056 17922 25057
rect 17606 24992 17612 25056
rect 17676 24992 17692 25056
rect 17756 24992 17772 25056
rect 17836 24992 17852 25056
rect 17916 24992 17922 25056
rect 17606 24991 17922 24992
rect 22606 25056 22922 25057
rect 22606 24992 22612 25056
rect 22676 24992 22692 25056
rect 22756 24992 22772 25056
rect 22836 24992 22852 25056
rect 22916 24992 22922 25056
rect 22606 24991 22922 24992
rect 27606 25056 27922 25057
rect 27606 24992 27612 25056
rect 27676 24992 27692 25056
rect 27756 24992 27772 25056
rect 27836 24992 27852 25056
rect 27916 24992 27922 25056
rect 27606 24991 27922 24992
rect 32606 25056 32922 25057
rect 32606 24992 32612 25056
rect 32676 24992 32692 25056
rect 32756 24992 32772 25056
rect 32836 24992 32852 25056
rect 32916 24992 32922 25056
rect 32606 24991 32922 24992
rect 37606 25056 37922 25057
rect 37606 24992 37612 25056
rect 37676 24992 37692 25056
rect 37756 24992 37772 25056
rect 37836 24992 37852 25056
rect 37916 24992 37922 25056
rect 37606 24991 37922 24992
rect 1946 24512 2262 24513
rect 1946 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2262 24512
rect 1946 24447 2262 24448
rect 6946 24512 7262 24513
rect 6946 24448 6952 24512
rect 7016 24448 7032 24512
rect 7096 24448 7112 24512
rect 7176 24448 7192 24512
rect 7256 24448 7262 24512
rect 6946 24447 7262 24448
rect 11946 24512 12262 24513
rect 11946 24448 11952 24512
rect 12016 24448 12032 24512
rect 12096 24448 12112 24512
rect 12176 24448 12192 24512
rect 12256 24448 12262 24512
rect 11946 24447 12262 24448
rect 16946 24512 17262 24513
rect 16946 24448 16952 24512
rect 17016 24448 17032 24512
rect 17096 24448 17112 24512
rect 17176 24448 17192 24512
rect 17256 24448 17262 24512
rect 16946 24447 17262 24448
rect 21946 24512 22262 24513
rect 21946 24448 21952 24512
rect 22016 24448 22032 24512
rect 22096 24448 22112 24512
rect 22176 24448 22192 24512
rect 22256 24448 22262 24512
rect 21946 24447 22262 24448
rect 26946 24512 27262 24513
rect 26946 24448 26952 24512
rect 27016 24448 27032 24512
rect 27096 24448 27112 24512
rect 27176 24448 27192 24512
rect 27256 24448 27262 24512
rect 26946 24447 27262 24448
rect 31946 24512 32262 24513
rect 31946 24448 31952 24512
rect 32016 24448 32032 24512
rect 32096 24448 32112 24512
rect 32176 24448 32192 24512
rect 32256 24448 32262 24512
rect 31946 24447 32262 24448
rect 36946 24512 37262 24513
rect 36946 24448 36952 24512
rect 37016 24448 37032 24512
rect 37096 24448 37112 24512
rect 37176 24448 37192 24512
rect 37256 24448 37262 24512
rect 36946 24447 37262 24448
rect 2606 23968 2922 23969
rect 2606 23904 2612 23968
rect 2676 23904 2692 23968
rect 2756 23904 2772 23968
rect 2836 23904 2852 23968
rect 2916 23904 2922 23968
rect 2606 23903 2922 23904
rect 7606 23968 7922 23969
rect 7606 23904 7612 23968
rect 7676 23904 7692 23968
rect 7756 23904 7772 23968
rect 7836 23904 7852 23968
rect 7916 23904 7922 23968
rect 7606 23903 7922 23904
rect 12606 23968 12922 23969
rect 12606 23904 12612 23968
rect 12676 23904 12692 23968
rect 12756 23904 12772 23968
rect 12836 23904 12852 23968
rect 12916 23904 12922 23968
rect 12606 23903 12922 23904
rect 17606 23968 17922 23969
rect 17606 23904 17612 23968
rect 17676 23904 17692 23968
rect 17756 23904 17772 23968
rect 17836 23904 17852 23968
rect 17916 23904 17922 23968
rect 17606 23903 17922 23904
rect 22606 23968 22922 23969
rect 22606 23904 22612 23968
rect 22676 23904 22692 23968
rect 22756 23904 22772 23968
rect 22836 23904 22852 23968
rect 22916 23904 22922 23968
rect 22606 23903 22922 23904
rect 27606 23968 27922 23969
rect 27606 23904 27612 23968
rect 27676 23904 27692 23968
rect 27756 23904 27772 23968
rect 27836 23904 27852 23968
rect 27916 23904 27922 23968
rect 27606 23903 27922 23904
rect 32606 23968 32922 23969
rect 32606 23904 32612 23968
rect 32676 23904 32692 23968
rect 32756 23904 32772 23968
rect 32836 23904 32852 23968
rect 32916 23904 32922 23968
rect 32606 23903 32922 23904
rect 37606 23968 37922 23969
rect 37606 23904 37612 23968
rect 37676 23904 37692 23968
rect 37756 23904 37772 23968
rect 37836 23904 37852 23968
rect 37916 23904 37922 23968
rect 37606 23903 37922 23904
rect 1946 23424 2262 23425
rect 1946 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2262 23424
rect 1946 23359 2262 23360
rect 6946 23424 7262 23425
rect 6946 23360 6952 23424
rect 7016 23360 7032 23424
rect 7096 23360 7112 23424
rect 7176 23360 7192 23424
rect 7256 23360 7262 23424
rect 6946 23359 7262 23360
rect 11946 23424 12262 23425
rect 11946 23360 11952 23424
rect 12016 23360 12032 23424
rect 12096 23360 12112 23424
rect 12176 23360 12192 23424
rect 12256 23360 12262 23424
rect 11946 23359 12262 23360
rect 16946 23424 17262 23425
rect 16946 23360 16952 23424
rect 17016 23360 17032 23424
rect 17096 23360 17112 23424
rect 17176 23360 17192 23424
rect 17256 23360 17262 23424
rect 16946 23359 17262 23360
rect 21946 23424 22262 23425
rect 21946 23360 21952 23424
rect 22016 23360 22032 23424
rect 22096 23360 22112 23424
rect 22176 23360 22192 23424
rect 22256 23360 22262 23424
rect 21946 23359 22262 23360
rect 26946 23424 27262 23425
rect 26946 23360 26952 23424
rect 27016 23360 27032 23424
rect 27096 23360 27112 23424
rect 27176 23360 27192 23424
rect 27256 23360 27262 23424
rect 26946 23359 27262 23360
rect 31946 23424 32262 23425
rect 31946 23360 31952 23424
rect 32016 23360 32032 23424
rect 32096 23360 32112 23424
rect 32176 23360 32192 23424
rect 32256 23360 32262 23424
rect 31946 23359 32262 23360
rect 36946 23424 37262 23425
rect 36946 23360 36952 23424
rect 37016 23360 37032 23424
rect 37096 23360 37112 23424
rect 37176 23360 37192 23424
rect 37256 23360 37262 23424
rect 36946 23359 37262 23360
rect 2606 22880 2922 22881
rect 2606 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2922 22880
rect 2606 22815 2922 22816
rect 7606 22880 7922 22881
rect 7606 22816 7612 22880
rect 7676 22816 7692 22880
rect 7756 22816 7772 22880
rect 7836 22816 7852 22880
rect 7916 22816 7922 22880
rect 7606 22815 7922 22816
rect 12606 22880 12922 22881
rect 12606 22816 12612 22880
rect 12676 22816 12692 22880
rect 12756 22816 12772 22880
rect 12836 22816 12852 22880
rect 12916 22816 12922 22880
rect 12606 22815 12922 22816
rect 17606 22880 17922 22881
rect 17606 22816 17612 22880
rect 17676 22816 17692 22880
rect 17756 22816 17772 22880
rect 17836 22816 17852 22880
rect 17916 22816 17922 22880
rect 17606 22815 17922 22816
rect 22606 22880 22922 22881
rect 22606 22816 22612 22880
rect 22676 22816 22692 22880
rect 22756 22816 22772 22880
rect 22836 22816 22852 22880
rect 22916 22816 22922 22880
rect 22606 22815 22922 22816
rect 27606 22880 27922 22881
rect 27606 22816 27612 22880
rect 27676 22816 27692 22880
rect 27756 22816 27772 22880
rect 27836 22816 27852 22880
rect 27916 22816 27922 22880
rect 27606 22815 27922 22816
rect 32606 22880 32922 22881
rect 32606 22816 32612 22880
rect 32676 22816 32692 22880
rect 32756 22816 32772 22880
rect 32836 22816 32852 22880
rect 32916 22816 32922 22880
rect 32606 22815 32922 22816
rect 37606 22880 37922 22881
rect 37606 22816 37612 22880
rect 37676 22816 37692 22880
rect 37756 22816 37772 22880
rect 37836 22816 37852 22880
rect 37916 22816 37922 22880
rect 37606 22815 37922 22816
rect 1946 22336 2262 22337
rect 1946 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2262 22336
rect 1946 22271 2262 22272
rect 6946 22336 7262 22337
rect 6946 22272 6952 22336
rect 7016 22272 7032 22336
rect 7096 22272 7112 22336
rect 7176 22272 7192 22336
rect 7256 22272 7262 22336
rect 6946 22271 7262 22272
rect 11946 22336 12262 22337
rect 11946 22272 11952 22336
rect 12016 22272 12032 22336
rect 12096 22272 12112 22336
rect 12176 22272 12192 22336
rect 12256 22272 12262 22336
rect 11946 22271 12262 22272
rect 16946 22336 17262 22337
rect 16946 22272 16952 22336
rect 17016 22272 17032 22336
rect 17096 22272 17112 22336
rect 17176 22272 17192 22336
rect 17256 22272 17262 22336
rect 16946 22271 17262 22272
rect 21946 22336 22262 22337
rect 21946 22272 21952 22336
rect 22016 22272 22032 22336
rect 22096 22272 22112 22336
rect 22176 22272 22192 22336
rect 22256 22272 22262 22336
rect 21946 22271 22262 22272
rect 26946 22336 27262 22337
rect 26946 22272 26952 22336
rect 27016 22272 27032 22336
rect 27096 22272 27112 22336
rect 27176 22272 27192 22336
rect 27256 22272 27262 22336
rect 26946 22271 27262 22272
rect 31946 22336 32262 22337
rect 31946 22272 31952 22336
rect 32016 22272 32032 22336
rect 32096 22272 32112 22336
rect 32176 22272 32192 22336
rect 32256 22272 32262 22336
rect 31946 22271 32262 22272
rect 36946 22336 37262 22337
rect 36946 22272 36952 22336
rect 37016 22272 37032 22336
rect 37096 22272 37112 22336
rect 37176 22272 37192 22336
rect 37256 22272 37262 22336
rect 36946 22271 37262 22272
rect 38469 21858 38535 21861
rect 39200 21858 40000 21888
rect 38469 21856 40000 21858
rect 38469 21800 38474 21856
rect 38530 21800 40000 21856
rect 38469 21798 40000 21800
rect 38469 21795 38535 21798
rect 2606 21792 2922 21793
rect 2606 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2922 21792
rect 2606 21727 2922 21728
rect 7606 21792 7922 21793
rect 7606 21728 7612 21792
rect 7676 21728 7692 21792
rect 7756 21728 7772 21792
rect 7836 21728 7852 21792
rect 7916 21728 7922 21792
rect 7606 21727 7922 21728
rect 12606 21792 12922 21793
rect 12606 21728 12612 21792
rect 12676 21728 12692 21792
rect 12756 21728 12772 21792
rect 12836 21728 12852 21792
rect 12916 21728 12922 21792
rect 12606 21727 12922 21728
rect 17606 21792 17922 21793
rect 17606 21728 17612 21792
rect 17676 21728 17692 21792
rect 17756 21728 17772 21792
rect 17836 21728 17852 21792
rect 17916 21728 17922 21792
rect 17606 21727 17922 21728
rect 22606 21792 22922 21793
rect 22606 21728 22612 21792
rect 22676 21728 22692 21792
rect 22756 21728 22772 21792
rect 22836 21728 22852 21792
rect 22916 21728 22922 21792
rect 22606 21727 22922 21728
rect 27606 21792 27922 21793
rect 27606 21728 27612 21792
rect 27676 21728 27692 21792
rect 27756 21728 27772 21792
rect 27836 21728 27852 21792
rect 27916 21728 27922 21792
rect 27606 21727 27922 21728
rect 32606 21792 32922 21793
rect 32606 21728 32612 21792
rect 32676 21728 32692 21792
rect 32756 21728 32772 21792
rect 32836 21728 32852 21792
rect 32916 21728 32922 21792
rect 32606 21727 32922 21728
rect 37606 21792 37922 21793
rect 37606 21728 37612 21792
rect 37676 21728 37692 21792
rect 37756 21728 37772 21792
rect 37836 21728 37852 21792
rect 37916 21728 37922 21792
rect 39200 21768 40000 21798
rect 37606 21727 37922 21728
rect 1946 21248 2262 21249
rect 0 21178 800 21208
rect 1946 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2262 21248
rect 1946 21183 2262 21184
rect 6946 21248 7262 21249
rect 6946 21184 6952 21248
rect 7016 21184 7032 21248
rect 7096 21184 7112 21248
rect 7176 21184 7192 21248
rect 7256 21184 7262 21248
rect 6946 21183 7262 21184
rect 11946 21248 12262 21249
rect 11946 21184 11952 21248
rect 12016 21184 12032 21248
rect 12096 21184 12112 21248
rect 12176 21184 12192 21248
rect 12256 21184 12262 21248
rect 11946 21183 12262 21184
rect 16946 21248 17262 21249
rect 16946 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17262 21248
rect 16946 21183 17262 21184
rect 21946 21248 22262 21249
rect 21946 21184 21952 21248
rect 22016 21184 22032 21248
rect 22096 21184 22112 21248
rect 22176 21184 22192 21248
rect 22256 21184 22262 21248
rect 21946 21183 22262 21184
rect 26946 21248 27262 21249
rect 26946 21184 26952 21248
rect 27016 21184 27032 21248
rect 27096 21184 27112 21248
rect 27176 21184 27192 21248
rect 27256 21184 27262 21248
rect 26946 21183 27262 21184
rect 31946 21248 32262 21249
rect 31946 21184 31952 21248
rect 32016 21184 32032 21248
rect 32096 21184 32112 21248
rect 32176 21184 32192 21248
rect 32256 21184 32262 21248
rect 31946 21183 32262 21184
rect 36946 21248 37262 21249
rect 36946 21184 36952 21248
rect 37016 21184 37032 21248
rect 37096 21184 37112 21248
rect 37176 21184 37192 21248
rect 37256 21184 37262 21248
rect 36946 21183 37262 21184
rect 933 21178 999 21181
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 38469 21178 38535 21181
rect 39200 21178 40000 21208
rect 38469 21176 40000 21178
rect 38469 21120 38474 21176
rect 38530 21120 40000 21176
rect 38469 21118 40000 21120
rect 38469 21115 38535 21118
rect 39200 21088 40000 21118
rect 2606 20704 2922 20705
rect 2606 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2922 20704
rect 2606 20639 2922 20640
rect 7606 20704 7922 20705
rect 7606 20640 7612 20704
rect 7676 20640 7692 20704
rect 7756 20640 7772 20704
rect 7836 20640 7852 20704
rect 7916 20640 7922 20704
rect 7606 20639 7922 20640
rect 12606 20704 12922 20705
rect 12606 20640 12612 20704
rect 12676 20640 12692 20704
rect 12756 20640 12772 20704
rect 12836 20640 12852 20704
rect 12916 20640 12922 20704
rect 12606 20639 12922 20640
rect 17606 20704 17922 20705
rect 17606 20640 17612 20704
rect 17676 20640 17692 20704
rect 17756 20640 17772 20704
rect 17836 20640 17852 20704
rect 17916 20640 17922 20704
rect 17606 20639 17922 20640
rect 22606 20704 22922 20705
rect 22606 20640 22612 20704
rect 22676 20640 22692 20704
rect 22756 20640 22772 20704
rect 22836 20640 22852 20704
rect 22916 20640 22922 20704
rect 22606 20639 22922 20640
rect 27606 20704 27922 20705
rect 27606 20640 27612 20704
rect 27676 20640 27692 20704
rect 27756 20640 27772 20704
rect 27836 20640 27852 20704
rect 27916 20640 27922 20704
rect 27606 20639 27922 20640
rect 32606 20704 32922 20705
rect 32606 20640 32612 20704
rect 32676 20640 32692 20704
rect 32756 20640 32772 20704
rect 32836 20640 32852 20704
rect 32916 20640 32922 20704
rect 32606 20639 32922 20640
rect 37606 20704 37922 20705
rect 37606 20640 37612 20704
rect 37676 20640 37692 20704
rect 37756 20640 37772 20704
rect 37836 20640 37852 20704
rect 37916 20640 37922 20704
rect 37606 20639 37922 20640
rect 1393 20634 1459 20637
rect 798 20632 1459 20634
rect 798 20576 1398 20632
rect 1454 20576 1459 20632
rect 798 20574 1459 20576
rect 798 20528 858 20574
rect 1393 20571 1459 20574
rect 0 20438 858 20528
rect 39021 20498 39087 20501
rect 39200 20498 40000 20528
rect 39021 20496 40000 20498
rect 39021 20440 39026 20496
rect 39082 20440 40000 20496
rect 39021 20438 40000 20440
rect 0 20408 800 20438
rect 39021 20435 39087 20438
rect 39200 20408 40000 20438
rect 1946 20160 2262 20161
rect 1946 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2262 20160
rect 1946 20095 2262 20096
rect 6946 20160 7262 20161
rect 6946 20096 6952 20160
rect 7016 20096 7032 20160
rect 7096 20096 7112 20160
rect 7176 20096 7192 20160
rect 7256 20096 7262 20160
rect 6946 20095 7262 20096
rect 11946 20160 12262 20161
rect 11946 20096 11952 20160
rect 12016 20096 12032 20160
rect 12096 20096 12112 20160
rect 12176 20096 12192 20160
rect 12256 20096 12262 20160
rect 11946 20095 12262 20096
rect 16946 20160 17262 20161
rect 16946 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17262 20160
rect 16946 20095 17262 20096
rect 21946 20160 22262 20161
rect 21946 20096 21952 20160
rect 22016 20096 22032 20160
rect 22096 20096 22112 20160
rect 22176 20096 22192 20160
rect 22256 20096 22262 20160
rect 21946 20095 22262 20096
rect 26946 20160 27262 20161
rect 26946 20096 26952 20160
rect 27016 20096 27032 20160
rect 27096 20096 27112 20160
rect 27176 20096 27192 20160
rect 27256 20096 27262 20160
rect 26946 20095 27262 20096
rect 31946 20160 32262 20161
rect 31946 20096 31952 20160
rect 32016 20096 32032 20160
rect 32096 20096 32112 20160
rect 32176 20096 32192 20160
rect 32256 20096 32262 20160
rect 31946 20095 32262 20096
rect 36946 20160 37262 20161
rect 36946 20096 36952 20160
rect 37016 20096 37032 20160
rect 37096 20096 37112 20160
rect 37176 20096 37192 20160
rect 37256 20096 37262 20160
rect 36946 20095 37262 20096
rect 0 19818 800 19848
rect 933 19818 999 19821
rect 0 19816 999 19818
rect 0 19760 938 19816
rect 994 19760 999 19816
rect 0 19758 999 19760
rect 0 19728 800 19758
rect 933 19755 999 19758
rect 38837 19818 38903 19821
rect 39200 19818 40000 19848
rect 38837 19816 40000 19818
rect 38837 19760 38842 19816
rect 38898 19760 40000 19816
rect 38837 19758 40000 19760
rect 38837 19755 38903 19758
rect 39200 19728 40000 19758
rect 2606 19616 2922 19617
rect 2606 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2922 19616
rect 2606 19551 2922 19552
rect 7606 19616 7922 19617
rect 7606 19552 7612 19616
rect 7676 19552 7692 19616
rect 7756 19552 7772 19616
rect 7836 19552 7852 19616
rect 7916 19552 7922 19616
rect 7606 19551 7922 19552
rect 12606 19616 12922 19617
rect 12606 19552 12612 19616
rect 12676 19552 12692 19616
rect 12756 19552 12772 19616
rect 12836 19552 12852 19616
rect 12916 19552 12922 19616
rect 12606 19551 12922 19552
rect 17606 19616 17922 19617
rect 17606 19552 17612 19616
rect 17676 19552 17692 19616
rect 17756 19552 17772 19616
rect 17836 19552 17852 19616
rect 17916 19552 17922 19616
rect 17606 19551 17922 19552
rect 22606 19616 22922 19617
rect 22606 19552 22612 19616
rect 22676 19552 22692 19616
rect 22756 19552 22772 19616
rect 22836 19552 22852 19616
rect 22916 19552 22922 19616
rect 22606 19551 22922 19552
rect 27606 19616 27922 19617
rect 27606 19552 27612 19616
rect 27676 19552 27692 19616
rect 27756 19552 27772 19616
rect 27836 19552 27852 19616
rect 27916 19552 27922 19616
rect 27606 19551 27922 19552
rect 32606 19616 32922 19617
rect 32606 19552 32612 19616
rect 32676 19552 32692 19616
rect 32756 19552 32772 19616
rect 32836 19552 32852 19616
rect 32916 19552 32922 19616
rect 32606 19551 32922 19552
rect 37606 19616 37922 19617
rect 37606 19552 37612 19616
rect 37676 19552 37692 19616
rect 37756 19552 37772 19616
rect 37836 19552 37852 19616
rect 37916 19552 37922 19616
rect 37606 19551 37922 19552
rect 18965 19410 19031 19413
rect 38285 19410 38351 19413
rect 18965 19408 38351 19410
rect 18965 19352 18970 19408
rect 19026 19352 38290 19408
rect 38346 19352 38351 19408
rect 18965 19350 38351 19352
rect 18965 19347 19031 19350
rect 38285 19347 38351 19350
rect 0 19138 800 19168
rect 1393 19138 1459 19141
rect 0 19136 1459 19138
rect 0 19080 1398 19136
rect 1454 19080 1459 19136
rect 0 19078 1459 19080
rect 0 19048 800 19078
rect 1393 19075 1459 19078
rect 38469 19138 38535 19141
rect 39200 19138 40000 19168
rect 38469 19136 40000 19138
rect 38469 19080 38474 19136
rect 38530 19080 40000 19136
rect 38469 19078 40000 19080
rect 38469 19075 38535 19078
rect 1946 19072 2262 19073
rect 1946 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2262 19072
rect 1946 19007 2262 19008
rect 6946 19072 7262 19073
rect 6946 19008 6952 19072
rect 7016 19008 7032 19072
rect 7096 19008 7112 19072
rect 7176 19008 7192 19072
rect 7256 19008 7262 19072
rect 6946 19007 7262 19008
rect 11946 19072 12262 19073
rect 11946 19008 11952 19072
rect 12016 19008 12032 19072
rect 12096 19008 12112 19072
rect 12176 19008 12192 19072
rect 12256 19008 12262 19072
rect 11946 19007 12262 19008
rect 16946 19072 17262 19073
rect 16946 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17262 19072
rect 16946 19007 17262 19008
rect 21946 19072 22262 19073
rect 21946 19008 21952 19072
rect 22016 19008 22032 19072
rect 22096 19008 22112 19072
rect 22176 19008 22192 19072
rect 22256 19008 22262 19072
rect 21946 19007 22262 19008
rect 26946 19072 27262 19073
rect 26946 19008 26952 19072
rect 27016 19008 27032 19072
rect 27096 19008 27112 19072
rect 27176 19008 27192 19072
rect 27256 19008 27262 19072
rect 26946 19007 27262 19008
rect 31946 19072 32262 19073
rect 31946 19008 31952 19072
rect 32016 19008 32032 19072
rect 32096 19008 32112 19072
rect 32176 19008 32192 19072
rect 32256 19008 32262 19072
rect 31946 19007 32262 19008
rect 36946 19072 37262 19073
rect 36946 19008 36952 19072
rect 37016 19008 37032 19072
rect 37096 19008 37112 19072
rect 37176 19008 37192 19072
rect 37256 19008 37262 19072
rect 39200 19048 40000 19078
rect 36946 19007 37262 19008
rect 2606 18528 2922 18529
rect 0 18458 800 18488
rect 2606 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2922 18528
rect 2606 18463 2922 18464
rect 7606 18528 7922 18529
rect 7606 18464 7612 18528
rect 7676 18464 7692 18528
rect 7756 18464 7772 18528
rect 7836 18464 7852 18528
rect 7916 18464 7922 18528
rect 7606 18463 7922 18464
rect 12606 18528 12922 18529
rect 12606 18464 12612 18528
rect 12676 18464 12692 18528
rect 12756 18464 12772 18528
rect 12836 18464 12852 18528
rect 12916 18464 12922 18528
rect 12606 18463 12922 18464
rect 17606 18528 17922 18529
rect 17606 18464 17612 18528
rect 17676 18464 17692 18528
rect 17756 18464 17772 18528
rect 17836 18464 17852 18528
rect 17916 18464 17922 18528
rect 17606 18463 17922 18464
rect 22606 18528 22922 18529
rect 22606 18464 22612 18528
rect 22676 18464 22692 18528
rect 22756 18464 22772 18528
rect 22836 18464 22852 18528
rect 22916 18464 22922 18528
rect 22606 18463 22922 18464
rect 27606 18528 27922 18529
rect 27606 18464 27612 18528
rect 27676 18464 27692 18528
rect 27756 18464 27772 18528
rect 27836 18464 27852 18528
rect 27916 18464 27922 18528
rect 27606 18463 27922 18464
rect 32606 18528 32922 18529
rect 32606 18464 32612 18528
rect 32676 18464 32692 18528
rect 32756 18464 32772 18528
rect 32836 18464 32852 18528
rect 32916 18464 32922 18528
rect 32606 18463 32922 18464
rect 37606 18528 37922 18529
rect 37606 18464 37612 18528
rect 37676 18464 37692 18528
rect 37756 18464 37772 18528
rect 37836 18464 37852 18528
rect 37916 18464 37922 18528
rect 37606 18463 37922 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 38469 18458 38535 18461
rect 39200 18458 40000 18488
rect 38469 18456 40000 18458
rect 38469 18400 38474 18456
rect 38530 18400 40000 18456
rect 38469 18398 40000 18400
rect 38469 18395 38535 18398
rect 39200 18368 40000 18398
rect 1946 17984 2262 17985
rect 1946 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2262 17984
rect 1946 17919 2262 17920
rect 6946 17984 7262 17985
rect 6946 17920 6952 17984
rect 7016 17920 7032 17984
rect 7096 17920 7112 17984
rect 7176 17920 7192 17984
rect 7256 17920 7262 17984
rect 6946 17919 7262 17920
rect 11946 17984 12262 17985
rect 11946 17920 11952 17984
rect 12016 17920 12032 17984
rect 12096 17920 12112 17984
rect 12176 17920 12192 17984
rect 12256 17920 12262 17984
rect 11946 17919 12262 17920
rect 16946 17984 17262 17985
rect 16946 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17262 17984
rect 16946 17919 17262 17920
rect 21946 17984 22262 17985
rect 21946 17920 21952 17984
rect 22016 17920 22032 17984
rect 22096 17920 22112 17984
rect 22176 17920 22192 17984
rect 22256 17920 22262 17984
rect 21946 17919 22262 17920
rect 26946 17984 27262 17985
rect 26946 17920 26952 17984
rect 27016 17920 27032 17984
rect 27096 17920 27112 17984
rect 27176 17920 27192 17984
rect 27256 17920 27262 17984
rect 26946 17919 27262 17920
rect 31946 17984 32262 17985
rect 31946 17920 31952 17984
rect 32016 17920 32032 17984
rect 32096 17920 32112 17984
rect 32176 17920 32192 17984
rect 32256 17920 32262 17984
rect 31946 17919 32262 17920
rect 36946 17984 37262 17985
rect 36946 17920 36952 17984
rect 37016 17920 37032 17984
rect 37096 17920 37112 17984
rect 37176 17920 37192 17984
rect 37256 17920 37262 17984
rect 36946 17919 37262 17920
rect 34513 17778 34579 17781
rect 39200 17778 40000 17808
rect 34513 17776 40000 17778
rect 34513 17720 34518 17776
rect 34574 17720 40000 17776
rect 34513 17718 40000 17720
rect 34513 17715 34579 17718
rect 39200 17688 40000 17718
rect 2606 17440 2922 17441
rect 2606 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2922 17440
rect 2606 17375 2922 17376
rect 7606 17440 7922 17441
rect 7606 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7922 17440
rect 7606 17375 7922 17376
rect 12606 17440 12922 17441
rect 12606 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12922 17440
rect 12606 17375 12922 17376
rect 17606 17440 17922 17441
rect 17606 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17922 17440
rect 17606 17375 17922 17376
rect 22606 17440 22922 17441
rect 22606 17376 22612 17440
rect 22676 17376 22692 17440
rect 22756 17376 22772 17440
rect 22836 17376 22852 17440
rect 22916 17376 22922 17440
rect 22606 17375 22922 17376
rect 27606 17440 27922 17441
rect 27606 17376 27612 17440
rect 27676 17376 27692 17440
rect 27756 17376 27772 17440
rect 27836 17376 27852 17440
rect 27916 17376 27922 17440
rect 27606 17375 27922 17376
rect 32606 17440 32922 17441
rect 32606 17376 32612 17440
rect 32676 17376 32692 17440
rect 32756 17376 32772 17440
rect 32836 17376 32852 17440
rect 32916 17376 32922 17440
rect 32606 17375 32922 17376
rect 37606 17440 37922 17441
rect 37606 17376 37612 17440
rect 37676 17376 37692 17440
rect 37756 17376 37772 17440
rect 37836 17376 37852 17440
rect 37916 17376 37922 17440
rect 37606 17375 37922 17376
rect 1946 16896 2262 16897
rect 1946 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2262 16896
rect 1946 16831 2262 16832
rect 6946 16896 7262 16897
rect 6946 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7262 16896
rect 6946 16831 7262 16832
rect 11946 16896 12262 16897
rect 11946 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12262 16896
rect 11946 16831 12262 16832
rect 16946 16896 17262 16897
rect 16946 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17262 16896
rect 16946 16831 17262 16832
rect 21946 16896 22262 16897
rect 21946 16832 21952 16896
rect 22016 16832 22032 16896
rect 22096 16832 22112 16896
rect 22176 16832 22192 16896
rect 22256 16832 22262 16896
rect 21946 16831 22262 16832
rect 26946 16896 27262 16897
rect 26946 16832 26952 16896
rect 27016 16832 27032 16896
rect 27096 16832 27112 16896
rect 27176 16832 27192 16896
rect 27256 16832 27262 16896
rect 26946 16831 27262 16832
rect 31946 16896 32262 16897
rect 31946 16832 31952 16896
rect 32016 16832 32032 16896
rect 32096 16832 32112 16896
rect 32176 16832 32192 16896
rect 32256 16832 32262 16896
rect 31946 16831 32262 16832
rect 36946 16896 37262 16897
rect 36946 16832 36952 16896
rect 37016 16832 37032 16896
rect 37096 16832 37112 16896
rect 37176 16832 37192 16896
rect 37256 16832 37262 16896
rect 36946 16831 37262 16832
rect 2606 16352 2922 16353
rect 2606 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2922 16352
rect 2606 16287 2922 16288
rect 7606 16352 7922 16353
rect 7606 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7922 16352
rect 7606 16287 7922 16288
rect 12606 16352 12922 16353
rect 12606 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12922 16352
rect 12606 16287 12922 16288
rect 17606 16352 17922 16353
rect 17606 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17922 16352
rect 17606 16287 17922 16288
rect 22606 16352 22922 16353
rect 22606 16288 22612 16352
rect 22676 16288 22692 16352
rect 22756 16288 22772 16352
rect 22836 16288 22852 16352
rect 22916 16288 22922 16352
rect 22606 16287 22922 16288
rect 27606 16352 27922 16353
rect 27606 16288 27612 16352
rect 27676 16288 27692 16352
rect 27756 16288 27772 16352
rect 27836 16288 27852 16352
rect 27916 16288 27922 16352
rect 27606 16287 27922 16288
rect 32606 16352 32922 16353
rect 32606 16288 32612 16352
rect 32676 16288 32692 16352
rect 32756 16288 32772 16352
rect 32836 16288 32852 16352
rect 32916 16288 32922 16352
rect 32606 16287 32922 16288
rect 37606 16352 37922 16353
rect 37606 16288 37612 16352
rect 37676 16288 37692 16352
rect 37756 16288 37772 16352
rect 37836 16288 37852 16352
rect 37916 16288 37922 16352
rect 37606 16287 37922 16288
rect 1946 15808 2262 15809
rect 1946 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2262 15808
rect 1946 15743 2262 15744
rect 6946 15808 7262 15809
rect 6946 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7262 15808
rect 6946 15743 7262 15744
rect 11946 15808 12262 15809
rect 11946 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12262 15808
rect 11946 15743 12262 15744
rect 16946 15808 17262 15809
rect 16946 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17262 15808
rect 16946 15743 17262 15744
rect 21946 15808 22262 15809
rect 21946 15744 21952 15808
rect 22016 15744 22032 15808
rect 22096 15744 22112 15808
rect 22176 15744 22192 15808
rect 22256 15744 22262 15808
rect 21946 15743 22262 15744
rect 26946 15808 27262 15809
rect 26946 15744 26952 15808
rect 27016 15744 27032 15808
rect 27096 15744 27112 15808
rect 27176 15744 27192 15808
rect 27256 15744 27262 15808
rect 26946 15743 27262 15744
rect 31946 15808 32262 15809
rect 31946 15744 31952 15808
rect 32016 15744 32032 15808
rect 32096 15744 32112 15808
rect 32176 15744 32192 15808
rect 32256 15744 32262 15808
rect 31946 15743 32262 15744
rect 36946 15808 37262 15809
rect 36946 15744 36952 15808
rect 37016 15744 37032 15808
rect 37096 15744 37112 15808
rect 37176 15744 37192 15808
rect 37256 15744 37262 15808
rect 36946 15743 37262 15744
rect 2606 15264 2922 15265
rect 2606 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2922 15264
rect 2606 15199 2922 15200
rect 7606 15264 7922 15265
rect 7606 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7922 15264
rect 7606 15199 7922 15200
rect 12606 15264 12922 15265
rect 12606 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12922 15264
rect 12606 15199 12922 15200
rect 17606 15264 17922 15265
rect 17606 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17922 15264
rect 17606 15199 17922 15200
rect 22606 15264 22922 15265
rect 22606 15200 22612 15264
rect 22676 15200 22692 15264
rect 22756 15200 22772 15264
rect 22836 15200 22852 15264
rect 22916 15200 22922 15264
rect 22606 15199 22922 15200
rect 27606 15264 27922 15265
rect 27606 15200 27612 15264
rect 27676 15200 27692 15264
rect 27756 15200 27772 15264
rect 27836 15200 27852 15264
rect 27916 15200 27922 15264
rect 27606 15199 27922 15200
rect 32606 15264 32922 15265
rect 32606 15200 32612 15264
rect 32676 15200 32692 15264
rect 32756 15200 32772 15264
rect 32836 15200 32852 15264
rect 32916 15200 32922 15264
rect 32606 15199 32922 15200
rect 37606 15264 37922 15265
rect 37606 15200 37612 15264
rect 37676 15200 37692 15264
rect 37756 15200 37772 15264
rect 37836 15200 37852 15264
rect 37916 15200 37922 15264
rect 37606 15199 37922 15200
rect 1946 14720 2262 14721
rect 1946 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2262 14720
rect 1946 14655 2262 14656
rect 6946 14720 7262 14721
rect 6946 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7262 14720
rect 6946 14655 7262 14656
rect 11946 14720 12262 14721
rect 11946 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12262 14720
rect 11946 14655 12262 14656
rect 16946 14720 17262 14721
rect 16946 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17262 14720
rect 16946 14655 17262 14656
rect 21946 14720 22262 14721
rect 21946 14656 21952 14720
rect 22016 14656 22032 14720
rect 22096 14656 22112 14720
rect 22176 14656 22192 14720
rect 22256 14656 22262 14720
rect 21946 14655 22262 14656
rect 26946 14720 27262 14721
rect 26946 14656 26952 14720
rect 27016 14656 27032 14720
rect 27096 14656 27112 14720
rect 27176 14656 27192 14720
rect 27256 14656 27262 14720
rect 26946 14655 27262 14656
rect 31946 14720 32262 14721
rect 31946 14656 31952 14720
rect 32016 14656 32032 14720
rect 32096 14656 32112 14720
rect 32176 14656 32192 14720
rect 32256 14656 32262 14720
rect 31946 14655 32262 14656
rect 36946 14720 37262 14721
rect 36946 14656 36952 14720
rect 37016 14656 37032 14720
rect 37096 14656 37112 14720
rect 37176 14656 37192 14720
rect 37256 14656 37262 14720
rect 36946 14655 37262 14656
rect 2606 14176 2922 14177
rect 2606 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2922 14176
rect 2606 14111 2922 14112
rect 7606 14176 7922 14177
rect 7606 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7922 14176
rect 7606 14111 7922 14112
rect 12606 14176 12922 14177
rect 12606 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12922 14176
rect 12606 14111 12922 14112
rect 17606 14176 17922 14177
rect 17606 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17922 14176
rect 17606 14111 17922 14112
rect 22606 14176 22922 14177
rect 22606 14112 22612 14176
rect 22676 14112 22692 14176
rect 22756 14112 22772 14176
rect 22836 14112 22852 14176
rect 22916 14112 22922 14176
rect 22606 14111 22922 14112
rect 27606 14176 27922 14177
rect 27606 14112 27612 14176
rect 27676 14112 27692 14176
rect 27756 14112 27772 14176
rect 27836 14112 27852 14176
rect 27916 14112 27922 14176
rect 27606 14111 27922 14112
rect 32606 14176 32922 14177
rect 32606 14112 32612 14176
rect 32676 14112 32692 14176
rect 32756 14112 32772 14176
rect 32836 14112 32852 14176
rect 32916 14112 32922 14176
rect 32606 14111 32922 14112
rect 37606 14176 37922 14177
rect 37606 14112 37612 14176
rect 37676 14112 37692 14176
rect 37756 14112 37772 14176
rect 37836 14112 37852 14176
rect 37916 14112 37922 14176
rect 37606 14111 37922 14112
rect 1946 13632 2262 13633
rect 1946 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2262 13632
rect 1946 13567 2262 13568
rect 6946 13632 7262 13633
rect 6946 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7262 13632
rect 6946 13567 7262 13568
rect 11946 13632 12262 13633
rect 11946 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12262 13632
rect 11946 13567 12262 13568
rect 16946 13632 17262 13633
rect 16946 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17262 13632
rect 16946 13567 17262 13568
rect 21946 13632 22262 13633
rect 21946 13568 21952 13632
rect 22016 13568 22032 13632
rect 22096 13568 22112 13632
rect 22176 13568 22192 13632
rect 22256 13568 22262 13632
rect 21946 13567 22262 13568
rect 26946 13632 27262 13633
rect 26946 13568 26952 13632
rect 27016 13568 27032 13632
rect 27096 13568 27112 13632
rect 27176 13568 27192 13632
rect 27256 13568 27262 13632
rect 26946 13567 27262 13568
rect 31946 13632 32262 13633
rect 31946 13568 31952 13632
rect 32016 13568 32032 13632
rect 32096 13568 32112 13632
rect 32176 13568 32192 13632
rect 32256 13568 32262 13632
rect 31946 13567 32262 13568
rect 36946 13632 37262 13633
rect 36946 13568 36952 13632
rect 37016 13568 37032 13632
rect 37096 13568 37112 13632
rect 37176 13568 37192 13632
rect 37256 13568 37262 13632
rect 36946 13567 37262 13568
rect 2606 13088 2922 13089
rect 2606 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2922 13088
rect 2606 13023 2922 13024
rect 7606 13088 7922 13089
rect 7606 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7922 13088
rect 7606 13023 7922 13024
rect 12606 13088 12922 13089
rect 12606 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12922 13088
rect 12606 13023 12922 13024
rect 17606 13088 17922 13089
rect 17606 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17922 13088
rect 17606 13023 17922 13024
rect 22606 13088 22922 13089
rect 22606 13024 22612 13088
rect 22676 13024 22692 13088
rect 22756 13024 22772 13088
rect 22836 13024 22852 13088
rect 22916 13024 22922 13088
rect 22606 13023 22922 13024
rect 27606 13088 27922 13089
rect 27606 13024 27612 13088
rect 27676 13024 27692 13088
rect 27756 13024 27772 13088
rect 27836 13024 27852 13088
rect 27916 13024 27922 13088
rect 27606 13023 27922 13024
rect 32606 13088 32922 13089
rect 32606 13024 32612 13088
rect 32676 13024 32692 13088
rect 32756 13024 32772 13088
rect 32836 13024 32852 13088
rect 32916 13024 32922 13088
rect 32606 13023 32922 13024
rect 37606 13088 37922 13089
rect 37606 13024 37612 13088
rect 37676 13024 37692 13088
rect 37756 13024 37772 13088
rect 37836 13024 37852 13088
rect 37916 13024 37922 13088
rect 37606 13023 37922 13024
rect 1946 12544 2262 12545
rect 1946 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2262 12544
rect 1946 12479 2262 12480
rect 6946 12544 7262 12545
rect 6946 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7262 12544
rect 6946 12479 7262 12480
rect 11946 12544 12262 12545
rect 11946 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12262 12544
rect 11946 12479 12262 12480
rect 16946 12544 17262 12545
rect 16946 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17262 12544
rect 16946 12479 17262 12480
rect 21946 12544 22262 12545
rect 21946 12480 21952 12544
rect 22016 12480 22032 12544
rect 22096 12480 22112 12544
rect 22176 12480 22192 12544
rect 22256 12480 22262 12544
rect 21946 12479 22262 12480
rect 26946 12544 27262 12545
rect 26946 12480 26952 12544
rect 27016 12480 27032 12544
rect 27096 12480 27112 12544
rect 27176 12480 27192 12544
rect 27256 12480 27262 12544
rect 26946 12479 27262 12480
rect 31946 12544 32262 12545
rect 31946 12480 31952 12544
rect 32016 12480 32032 12544
rect 32096 12480 32112 12544
rect 32176 12480 32192 12544
rect 32256 12480 32262 12544
rect 31946 12479 32262 12480
rect 36946 12544 37262 12545
rect 36946 12480 36952 12544
rect 37016 12480 37032 12544
rect 37096 12480 37112 12544
rect 37176 12480 37192 12544
rect 37256 12480 37262 12544
rect 36946 12479 37262 12480
rect 2606 12000 2922 12001
rect 2606 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2922 12000
rect 2606 11935 2922 11936
rect 7606 12000 7922 12001
rect 7606 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7922 12000
rect 7606 11935 7922 11936
rect 12606 12000 12922 12001
rect 12606 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12922 12000
rect 12606 11935 12922 11936
rect 17606 12000 17922 12001
rect 17606 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17922 12000
rect 17606 11935 17922 11936
rect 22606 12000 22922 12001
rect 22606 11936 22612 12000
rect 22676 11936 22692 12000
rect 22756 11936 22772 12000
rect 22836 11936 22852 12000
rect 22916 11936 22922 12000
rect 22606 11935 22922 11936
rect 27606 12000 27922 12001
rect 27606 11936 27612 12000
rect 27676 11936 27692 12000
rect 27756 11936 27772 12000
rect 27836 11936 27852 12000
rect 27916 11936 27922 12000
rect 27606 11935 27922 11936
rect 32606 12000 32922 12001
rect 32606 11936 32612 12000
rect 32676 11936 32692 12000
rect 32756 11936 32772 12000
rect 32836 11936 32852 12000
rect 32916 11936 32922 12000
rect 32606 11935 32922 11936
rect 37606 12000 37922 12001
rect 37606 11936 37612 12000
rect 37676 11936 37692 12000
rect 37756 11936 37772 12000
rect 37836 11936 37852 12000
rect 37916 11936 37922 12000
rect 37606 11935 37922 11936
rect 1946 11456 2262 11457
rect 1946 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2262 11456
rect 1946 11391 2262 11392
rect 6946 11456 7262 11457
rect 6946 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7262 11456
rect 6946 11391 7262 11392
rect 11946 11456 12262 11457
rect 11946 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12262 11456
rect 11946 11391 12262 11392
rect 16946 11456 17262 11457
rect 16946 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17262 11456
rect 16946 11391 17262 11392
rect 21946 11456 22262 11457
rect 21946 11392 21952 11456
rect 22016 11392 22032 11456
rect 22096 11392 22112 11456
rect 22176 11392 22192 11456
rect 22256 11392 22262 11456
rect 21946 11391 22262 11392
rect 26946 11456 27262 11457
rect 26946 11392 26952 11456
rect 27016 11392 27032 11456
rect 27096 11392 27112 11456
rect 27176 11392 27192 11456
rect 27256 11392 27262 11456
rect 26946 11391 27262 11392
rect 31946 11456 32262 11457
rect 31946 11392 31952 11456
rect 32016 11392 32032 11456
rect 32096 11392 32112 11456
rect 32176 11392 32192 11456
rect 32256 11392 32262 11456
rect 31946 11391 32262 11392
rect 36946 11456 37262 11457
rect 36946 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37262 11456
rect 36946 11391 37262 11392
rect 2606 10912 2922 10913
rect 2606 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2922 10912
rect 2606 10847 2922 10848
rect 7606 10912 7922 10913
rect 7606 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7922 10912
rect 7606 10847 7922 10848
rect 12606 10912 12922 10913
rect 12606 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12922 10912
rect 12606 10847 12922 10848
rect 17606 10912 17922 10913
rect 17606 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17922 10912
rect 17606 10847 17922 10848
rect 22606 10912 22922 10913
rect 22606 10848 22612 10912
rect 22676 10848 22692 10912
rect 22756 10848 22772 10912
rect 22836 10848 22852 10912
rect 22916 10848 22922 10912
rect 22606 10847 22922 10848
rect 27606 10912 27922 10913
rect 27606 10848 27612 10912
rect 27676 10848 27692 10912
rect 27756 10848 27772 10912
rect 27836 10848 27852 10912
rect 27916 10848 27922 10912
rect 27606 10847 27922 10848
rect 32606 10912 32922 10913
rect 32606 10848 32612 10912
rect 32676 10848 32692 10912
rect 32756 10848 32772 10912
rect 32836 10848 32852 10912
rect 32916 10848 32922 10912
rect 32606 10847 32922 10848
rect 37606 10912 37922 10913
rect 37606 10848 37612 10912
rect 37676 10848 37692 10912
rect 37756 10848 37772 10912
rect 37836 10848 37852 10912
rect 37916 10848 37922 10912
rect 37606 10847 37922 10848
rect 1946 10368 2262 10369
rect 1946 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2262 10368
rect 1946 10303 2262 10304
rect 6946 10368 7262 10369
rect 6946 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7262 10368
rect 6946 10303 7262 10304
rect 11946 10368 12262 10369
rect 11946 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12262 10368
rect 11946 10303 12262 10304
rect 16946 10368 17262 10369
rect 16946 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17262 10368
rect 16946 10303 17262 10304
rect 21946 10368 22262 10369
rect 21946 10304 21952 10368
rect 22016 10304 22032 10368
rect 22096 10304 22112 10368
rect 22176 10304 22192 10368
rect 22256 10304 22262 10368
rect 21946 10303 22262 10304
rect 26946 10368 27262 10369
rect 26946 10304 26952 10368
rect 27016 10304 27032 10368
rect 27096 10304 27112 10368
rect 27176 10304 27192 10368
rect 27256 10304 27262 10368
rect 26946 10303 27262 10304
rect 31946 10368 32262 10369
rect 31946 10304 31952 10368
rect 32016 10304 32032 10368
rect 32096 10304 32112 10368
rect 32176 10304 32192 10368
rect 32256 10304 32262 10368
rect 31946 10303 32262 10304
rect 36946 10368 37262 10369
rect 36946 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37262 10368
rect 36946 10303 37262 10304
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 7606 9824 7922 9825
rect 7606 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7922 9824
rect 7606 9759 7922 9760
rect 12606 9824 12922 9825
rect 12606 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12922 9824
rect 12606 9759 12922 9760
rect 17606 9824 17922 9825
rect 17606 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17922 9824
rect 17606 9759 17922 9760
rect 22606 9824 22922 9825
rect 22606 9760 22612 9824
rect 22676 9760 22692 9824
rect 22756 9760 22772 9824
rect 22836 9760 22852 9824
rect 22916 9760 22922 9824
rect 22606 9759 22922 9760
rect 27606 9824 27922 9825
rect 27606 9760 27612 9824
rect 27676 9760 27692 9824
rect 27756 9760 27772 9824
rect 27836 9760 27852 9824
rect 27916 9760 27922 9824
rect 27606 9759 27922 9760
rect 32606 9824 32922 9825
rect 32606 9760 32612 9824
rect 32676 9760 32692 9824
rect 32756 9760 32772 9824
rect 32836 9760 32852 9824
rect 32916 9760 32922 9824
rect 32606 9759 32922 9760
rect 37606 9824 37922 9825
rect 37606 9760 37612 9824
rect 37676 9760 37692 9824
rect 37756 9760 37772 9824
rect 37836 9760 37852 9824
rect 37916 9760 37922 9824
rect 37606 9759 37922 9760
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 6946 9280 7262 9281
rect 6946 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7262 9280
rect 6946 9215 7262 9216
rect 11946 9280 12262 9281
rect 11946 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12262 9280
rect 11946 9215 12262 9216
rect 16946 9280 17262 9281
rect 16946 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17262 9280
rect 16946 9215 17262 9216
rect 21946 9280 22262 9281
rect 21946 9216 21952 9280
rect 22016 9216 22032 9280
rect 22096 9216 22112 9280
rect 22176 9216 22192 9280
rect 22256 9216 22262 9280
rect 21946 9215 22262 9216
rect 26946 9280 27262 9281
rect 26946 9216 26952 9280
rect 27016 9216 27032 9280
rect 27096 9216 27112 9280
rect 27176 9216 27192 9280
rect 27256 9216 27262 9280
rect 26946 9215 27262 9216
rect 31946 9280 32262 9281
rect 31946 9216 31952 9280
rect 32016 9216 32032 9280
rect 32096 9216 32112 9280
rect 32176 9216 32192 9280
rect 32256 9216 32262 9280
rect 31946 9215 32262 9216
rect 36946 9280 37262 9281
rect 36946 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37262 9280
rect 36946 9215 37262 9216
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 7606 8736 7922 8737
rect 7606 8672 7612 8736
rect 7676 8672 7692 8736
rect 7756 8672 7772 8736
rect 7836 8672 7852 8736
rect 7916 8672 7922 8736
rect 7606 8671 7922 8672
rect 12606 8736 12922 8737
rect 12606 8672 12612 8736
rect 12676 8672 12692 8736
rect 12756 8672 12772 8736
rect 12836 8672 12852 8736
rect 12916 8672 12922 8736
rect 12606 8671 12922 8672
rect 17606 8736 17922 8737
rect 17606 8672 17612 8736
rect 17676 8672 17692 8736
rect 17756 8672 17772 8736
rect 17836 8672 17852 8736
rect 17916 8672 17922 8736
rect 17606 8671 17922 8672
rect 22606 8736 22922 8737
rect 22606 8672 22612 8736
rect 22676 8672 22692 8736
rect 22756 8672 22772 8736
rect 22836 8672 22852 8736
rect 22916 8672 22922 8736
rect 22606 8671 22922 8672
rect 27606 8736 27922 8737
rect 27606 8672 27612 8736
rect 27676 8672 27692 8736
rect 27756 8672 27772 8736
rect 27836 8672 27852 8736
rect 27916 8672 27922 8736
rect 27606 8671 27922 8672
rect 32606 8736 32922 8737
rect 32606 8672 32612 8736
rect 32676 8672 32692 8736
rect 32756 8672 32772 8736
rect 32836 8672 32852 8736
rect 32916 8672 32922 8736
rect 32606 8671 32922 8672
rect 37606 8736 37922 8737
rect 37606 8672 37612 8736
rect 37676 8672 37692 8736
rect 37756 8672 37772 8736
rect 37836 8672 37852 8736
rect 37916 8672 37922 8736
rect 37606 8671 37922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 6946 8192 7262 8193
rect 6946 8128 6952 8192
rect 7016 8128 7032 8192
rect 7096 8128 7112 8192
rect 7176 8128 7192 8192
rect 7256 8128 7262 8192
rect 6946 8127 7262 8128
rect 11946 8192 12262 8193
rect 11946 8128 11952 8192
rect 12016 8128 12032 8192
rect 12096 8128 12112 8192
rect 12176 8128 12192 8192
rect 12256 8128 12262 8192
rect 11946 8127 12262 8128
rect 16946 8192 17262 8193
rect 16946 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17262 8192
rect 16946 8127 17262 8128
rect 21946 8192 22262 8193
rect 21946 8128 21952 8192
rect 22016 8128 22032 8192
rect 22096 8128 22112 8192
rect 22176 8128 22192 8192
rect 22256 8128 22262 8192
rect 21946 8127 22262 8128
rect 26946 8192 27262 8193
rect 26946 8128 26952 8192
rect 27016 8128 27032 8192
rect 27096 8128 27112 8192
rect 27176 8128 27192 8192
rect 27256 8128 27262 8192
rect 26946 8127 27262 8128
rect 31946 8192 32262 8193
rect 31946 8128 31952 8192
rect 32016 8128 32032 8192
rect 32096 8128 32112 8192
rect 32176 8128 32192 8192
rect 32256 8128 32262 8192
rect 31946 8127 32262 8128
rect 36946 8192 37262 8193
rect 36946 8128 36952 8192
rect 37016 8128 37032 8192
rect 37096 8128 37112 8192
rect 37176 8128 37192 8192
rect 37256 8128 37262 8192
rect 36946 8127 37262 8128
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 7606 7648 7922 7649
rect 7606 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7922 7648
rect 7606 7583 7922 7584
rect 12606 7648 12922 7649
rect 12606 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12922 7648
rect 12606 7583 12922 7584
rect 17606 7648 17922 7649
rect 17606 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17922 7648
rect 17606 7583 17922 7584
rect 22606 7648 22922 7649
rect 22606 7584 22612 7648
rect 22676 7584 22692 7648
rect 22756 7584 22772 7648
rect 22836 7584 22852 7648
rect 22916 7584 22922 7648
rect 22606 7583 22922 7584
rect 27606 7648 27922 7649
rect 27606 7584 27612 7648
rect 27676 7584 27692 7648
rect 27756 7584 27772 7648
rect 27836 7584 27852 7648
rect 27916 7584 27922 7648
rect 27606 7583 27922 7584
rect 32606 7648 32922 7649
rect 32606 7584 32612 7648
rect 32676 7584 32692 7648
rect 32756 7584 32772 7648
rect 32836 7584 32852 7648
rect 32916 7584 32922 7648
rect 32606 7583 32922 7584
rect 37606 7648 37922 7649
rect 37606 7584 37612 7648
rect 37676 7584 37692 7648
rect 37756 7584 37772 7648
rect 37836 7584 37852 7648
rect 37916 7584 37922 7648
rect 37606 7583 37922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 6946 7104 7262 7105
rect 6946 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7262 7104
rect 6946 7039 7262 7040
rect 11946 7104 12262 7105
rect 11946 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12262 7104
rect 11946 7039 12262 7040
rect 16946 7104 17262 7105
rect 16946 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17262 7104
rect 16946 7039 17262 7040
rect 21946 7104 22262 7105
rect 21946 7040 21952 7104
rect 22016 7040 22032 7104
rect 22096 7040 22112 7104
rect 22176 7040 22192 7104
rect 22256 7040 22262 7104
rect 21946 7039 22262 7040
rect 26946 7104 27262 7105
rect 26946 7040 26952 7104
rect 27016 7040 27032 7104
rect 27096 7040 27112 7104
rect 27176 7040 27192 7104
rect 27256 7040 27262 7104
rect 26946 7039 27262 7040
rect 31946 7104 32262 7105
rect 31946 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32262 7104
rect 31946 7039 32262 7040
rect 36946 7104 37262 7105
rect 36946 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37262 7104
rect 36946 7039 37262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 7606 6560 7922 6561
rect 7606 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7922 6560
rect 7606 6495 7922 6496
rect 12606 6560 12922 6561
rect 12606 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12922 6560
rect 12606 6495 12922 6496
rect 17606 6560 17922 6561
rect 17606 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17922 6560
rect 17606 6495 17922 6496
rect 22606 6560 22922 6561
rect 22606 6496 22612 6560
rect 22676 6496 22692 6560
rect 22756 6496 22772 6560
rect 22836 6496 22852 6560
rect 22916 6496 22922 6560
rect 22606 6495 22922 6496
rect 27606 6560 27922 6561
rect 27606 6496 27612 6560
rect 27676 6496 27692 6560
rect 27756 6496 27772 6560
rect 27836 6496 27852 6560
rect 27916 6496 27922 6560
rect 27606 6495 27922 6496
rect 32606 6560 32922 6561
rect 32606 6496 32612 6560
rect 32676 6496 32692 6560
rect 32756 6496 32772 6560
rect 32836 6496 32852 6560
rect 32916 6496 32922 6560
rect 32606 6495 32922 6496
rect 37606 6560 37922 6561
rect 37606 6496 37612 6560
rect 37676 6496 37692 6560
rect 37756 6496 37772 6560
rect 37836 6496 37852 6560
rect 37916 6496 37922 6560
rect 37606 6495 37922 6496
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 6946 6016 7262 6017
rect 6946 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7262 6016
rect 6946 5951 7262 5952
rect 11946 6016 12262 6017
rect 11946 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12262 6016
rect 11946 5951 12262 5952
rect 16946 6016 17262 6017
rect 16946 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17262 6016
rect 16946 5951 17262 5952
rect 21946 6016 22262 6017
rect 21946 5952 21952 6016
rect 22016 5952 22032 6016
rect 22096 5952 22112 6016
rect 22176 5952 22192 6016
rect 22256 5952 22262 6016
rect 21946 5951 22262 5952
rect 26946 6016 27262 6017
rect 26946 5952 26952 6016
rect 27016 5952 27032 6016
rect 27096 5952 27112 6016
rect 27176 5952 27192 6016
rect 27256 5952 27262 6016
rect 26946 5951 27262 5952
rect 31946 6016 32262 6017
rect 31946 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32262 6016
rect 31946 5951 32262 5952
rect 36946 6016 37262 6017
rect 36946 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37262 6016
rect 36946 5951 37262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 7606 5472 7922 5473
rect 7606 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7922 5472
rect 7606 5407 7922 5408
rect 12606 5472 12922 5473
rect 12606 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12922 5472
rect 12606 5407 12922 5408
rect 17606 5472 17922 5473
rect 17606 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17922 5472
rect 17606 5407 17922 5408
rect 22606 5472 22922 5473
rect 22606 5408 22612 5472
rect 22676 5408 22692 5472
rect 22756 5408 22772 5472
rect 22836 5408 22852 5472
rect 22916 5408 22922 5472
rect 22606 5407 22922 5408
rect 27606 5472 27922 5473
rect 27606 5408 27612 5472
rect 27676 5408 27692 5472
rect 27756 5408 27772 5472
rect 27836 5408 27852 5472
rect 27916 5408 27922 5472
rect 27606 5407 27922 5408
rect 32606 5472 32922 5473
rect 32606 5408 32612 5472
rect 32676 5408 32692 5472
rect 32756 5408 32772 5472
rect 32836 5408 32852 5472
rect 32916 5408 32922 5472
rect 32606 5407 32922 5408
rect 37606 5472 37922 5473
rect 37606 5408 37612 5472
rect 37676 5408 37692 5472
rect 37756 5408 37772 5472
rect 37836 5408 37852 5472
rect 37916 5408 37922 5472
rect 37606 5407 37922 5408
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 6946 4928 7262 4929
rect 6946 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7262 4928
rect 6946 4863 7262 4864
rect 11946 4928 12262 4929
rect 11946 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12262 4928
rect 11946 4863 12262 4864
rect 16946 4928 17262 4929
rect 16946 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17262 4928
rect 16946 4863 17262 4864
rect 21946 4928 22262 4929
rect 21946 4864 21952 4928
rect 22016 4864 22032 4928
rect 22096 4864 22112 4928
rect 22176 4864 22192 4928
rect 22256 4864 22262 4928
rect 21946 4863 22262 4864
rect 26946 4928 27262 4929
rect 26946 4864 26952 4928
rect 27016 4864 27032 4928
rect 27096 4864 27112 4928
rect 27176 4864 27192 4928
rect 27256 4864 27262 4928
rect 26946 4863 27262 4864
rect 31946 4928 32262 4929
rect 31946 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32262 4928
rect 31946 4863 32262 4864
rect 36946 4928 37262 4929
rect 36946 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37262 4928
rect 36946 4863 37262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 7606 4384 7922 4385
rect 7606 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7922 4384
rect 7606 4319 7922 4320
rect 12606 4384 12922 4385
rect 12606 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12922 4384
rect 12606 4319 12922 4320
rect 17606 4384 17922 4385
rect 17606 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17922 4384
rect 17606 4319 17922 4320
rect 22606 4384 22922 4385
rect 22606 4320 22612 4384
rect 22676 4320 22692 4384
rect 22756 4320 22772 4384
rect 22836 4320 22852 4384
rect 22916 4320 22922 4384
rect 22606 4319 22922 4320
rect 27606 4384 27922 4385
rect 27606 4320 27612 4384
rect 27676 4320 27692 4384
rect 27756 4320 27772 4384
rect 27836 4320 27852 4384
rect 27916 4320 27922 4384
rect 27606 4319 27922 4320
rect 32606 4384 32922 4385
rect 32606 4320 32612 4384
rect 32676 4320 32692 4384
rect 32756 4320 32772 4384
rect 32836 4320 32852 4384
rect 32916 4320 32922 4384
rect 32606 4319 32922 4320
rect 37606 4384 37922 4385
rect 37606 4320 37612 4384
rect 37676 4320 37692 4384
rect 37756 4320 37772 4384
rect 37836 4320 37852 4384
rect 37916 4320 37922 4384
rect 37606 4319 37922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 6946 3840 7262 3841
rect 6946 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7262 3840
rect 6946 3775 7262 3776
rect 11946 3840 12262 3841
rect 11946 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12262 3840
rect 11946 3775 12262 3776
rect 16946 3840 17262 3841
rect 16946 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17262 3840
rect 16946 3775 17262 3776
rect 21946 3840 22262 3841
rect 21946 3776 21952 3840
rect 22016 3776 22032 3840
rect 22096 3776 22112 3840
rect 22176 3776 22192 3840
rect 22256 3776 22262 3840
rect 21946 3775 22262 3776
rect 26946 3840 27262 3841
rect 26946 3776 26952 3840
rect 27016 3776 27032 3840
rect 27096 3776 27112 3840
rect 27176 3776 27192 3840
rect 27256 3776 27262 3840
rect 26946 3775 27262 3776
rect 31946 3840 32262 3841
rect 31946 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32262 3840
rect 31946 3775 32262 3776
rect 36946 3840 37262 3841
rect 36946 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37262 3840
rect 36946 3775 37262 3776
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 7606 3296 7922 3297
rect 7606 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7922 3296
rect 7606 3231 7922 3232
rect 12606 3296 12922 3297
rect 12606 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12922 3296
rect 12606 3231 12922 3232
rect 17606 3296 17922 3297
rect 17606 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17922 3296
rect 17606 3231 17922 3232
rect 22606 3296 22922 3297
rect 22606 3232 22612 3296
rect 22676 3232 22692 3296
rect 22756 3232 22772 3296
rect 22836 3232 22852 3296
rect 22916 3232 22922 3296
rect 22606 3231 22922 3232
rect 27606 3296 27922 3297
rect 27606 3232 27612 3296
rect 27676 3232 27692 3296
rect 27756 3232 27772 3296
rect 27836 3232 27852 3296
rect 27916 3232 27922 3296
rect 27606 3231 27922 3232
rect 32606 3296 32922 3297
rect 32606 3232 32612 3296
rect 32676 3232 32692 3296
rect 32756 3232 32772 3296
rect 32836 3232 32852 3296
rect 32916 3232 32922 3296
rect 32606 3231 32922 3232
rect 37606 3296 37922 3297
rect 37606 3232 37612 3296
rect 37676 3232 37692 3296
rect 37756 3232 37772 3296
rect 37836 3232 37852 3296
rect 37916 3232 37922 3296
rect 37606 3231 37922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 6946 2752 7262 2753
rect 6946 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7262 2752
rect 6946 2687 7262 2688
rect 11946 2752 12262 2753
rect 11946 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12262 2752
rect 11946 2687 12262 2688
rect 16946 2752 17262 2753
rect 16946 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17262 2752
rect 16946 2687 17262 2688
rect 21946 2752 22262 2753
rect 21946 2688 21952 2752
rect 22016 2688 22032 2752
rect 22096 2688 22112 2752
rect 22176 2688 22192 2752
rect 22256 2688 22262 2752
rect 21946 2687 22262 2688
rect 26946 2752 27262 2753
rect 26946 2688 26952 2752
rect 27016 2688 27032 2752
rect 27096 2688 27112 2752
rect 27176 2688 27192 2752
rect 27256 2688 27262 2752
rect 26946 2687 27262 2688
rect 31946 2752 32262 2753
rect 31946 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32262 2752
rect 31946 2687 32262 2688
rect 36946 2752 37262 2753
rect 36946 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37262 2752
rect 36946 2687 37262 2688
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 7606 2208 7922 2209
rect 7606 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7922 2208
rect 7606 2143 7922 2144
rect 12606 2208 12922 2209
rect 12606 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12922 2208
rect 12606 2143 12922 2144
rect 17606 2208 17922 2209
rect 17606 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17922 2208
rect 17606 2143 17922 2144
rect 22606 2208 22922 2209
rect 22606 2144 22612 2208
rect 22676 2144 22692 2208
rect 22756 2144 22772 2208
rect 22836 2144 22852 2208
rect 22916 2144 22922 2208
rect 22606 2143 22922 2144
rect 27606 2208 27922 2209
rect 27606 2144 27612 2208
rect 27676 2144 27692 2208
rect 27756 2144 27772 2208
rect 27836 2144 27852 2208
rect 27916 2144 27922 2208
rect 27606 2143 27922 2144
rect 32606 2208 32922 2209
rect 32606 2144 32612 2208
rect 32676 2144 32692 2208
rect 32756 2144 32772 2208
rect 32836 2144 32852 2208
rect 32916 2144 32922 2208
rect 32606 2143 32922 2144
rect 37606 2208 37922 2209
rect 37606 2144 37612 2208
rect 37676 2144 37692 2208
rect 37756 2144 37772 2208
rect 37836 2144 37852 2208
rect 37916 2144 37922 2208
rect 37606 2143 37922 2144
<< via3 >>
rect 1952 37564 2016 37568
rect 1952 37508 1956 37564
rect 1956 37508 2012 37564
rect 2012 37508 2016 37564
rect 1952 37504 2016 37508
rect 2032 37564 2096 37568
rect 2032 37508 2036 37564
rect 2036 37508 2092 37564
rect 2092 37508 2096 37564
rect 2032 37504 2096 37508
rect 2112 37564 2176 37568
rect 2112 37508 2116 37564
rect 2116 37508 2172 37564
rect 2172 37508 2176 37564
rect 2112 37504 2176 37508
rect 2192 37564 2256 37568
rect 2192 37508 2196 37564
rect 2196 37508 2252 37564
rect 2252 37508 2256 37564
rect 2192 37504 2256 37508
rect 6952 37564 7016 37568
rect 6952 37508 6956 37564
rect 6956 37508 7012 37564
rect 7012 37508 7016 37564
rect 6952 37504 7016 37508
rect 7032 37564 7096 37568
rect 7032 37508 7036 37564
rect 7036 37508 7092 37564
rect 7092 37508 7096 37564
rect 7032 37504 7096 37508
rect 7112 37564 7176 37568
rect 7112 37508 7116 37564
rect 7116 37508 7172 37564
rect 7172 37508 7176 37564
rect 7112 37504 7176 37508
rect 7192 37564 7256 37568
rect 7192 37508 7196 37564
rect 7196 37508 7252 37564
rect 7252 37508 7256 37564
rect 7192 37504 7256 37508
rect 11952 37564 12016 37568
rect 11952 37508 11956 37564
rect 11956 37508 12012 37564
rect 12012 37508 12016 37564
rect 11952 37504 12016 37508
rect 12032 37564 12096 37568
rect 12032 37508 12036 37564
rect 12036 37508 12092 37564
rect 12092 37508 12096 37564
rect 12032 37504 12096 37508
rect 12112 37564 12176 37568
rect 12112 37508 12116 37564
rect 12116 37508 12172 37564
rect 12172 37508 12176 37564
rect 12112 37504 12176 37508
rect 12192 37564 12256 37568
rect 12192 37508 12196 37564
rect 12196 37508 12252 37564
rect 12252 37508 12256 37564
rect 12192 37504 12256 37508
rect 16952 37564 17016 37568
rect 16952 37508 16956 37564
rect 16956 37508 17012 37564
rect 17012 37508 17016 37564
rect 16952 37504 17016 37508
rect 17032 37564 17096 37568
rect 17032 37508 17036 37564
rect 17036 37508 17092 37564
rect 17092 37508 17096 37564
rect 17032 37504 17096 37508
rect 17112 37564 17176 37568
rect 17112 37508 17116 37564
rect 17116 37508 17172 37564
rect 17172 37508 17176 37564
rect 17112 37504 17176 37508
rect 17192 37564 17256 37568
rect 17192 37508 17196 37564
rect 17196 37508 17252 37564
rect 17252 37508 17256 37564
rect 17192 37504 17256 37508
rect 21952 37564 22016 37568
rect 21952 37508 21956 37564
rect 21956 37508 22012 37564
rect 22012 37508 22016 37564
rect 21952 37504 22016 37508
rect 22032 37564 22096 37568
rect 22032 37508 22036 37564
rect 22036 37508 22092 37564
rect 22092 37508 22096 37564
rect 22032 37504 22096 37508
rect 22112 37564 22176 37568
rect 22112 37508 22116 37564
rect 22116 37508 22172 37564
rect 22172 37508 22176 37564
rect 22112 37504 22176 37508
rect 22192 37564 22256 37568
rect 22192 37508 22196 37564
rect 22196 37508 22252 37564
rect 22252 37508 22256 37564
rect 22192 37504 22256 37508
rect 26952 37564 27016 37568
rect 26952 37508 26956 37564
rect 26956 37508 27012 37564
rect 27012 37508 27016 37564
rect 26952 37504 27016 37508
rect 27032 37564 27096 37568
rect 27032 37508 27036 37564
rect 27036 37508 27092 37564
rect 27092 37508 27096 37564
rect 27032 37504 27096 37508
rect 27112 37564 27176 37568
rect 27112 37508 27116 37564
rect 27116 37508 27172 37564
rect 27172 37508 27176 37564
rect 27112 37504 27176 37508
rect 27192 37564 27256 37568
rect 27192 37508 27196 37564
rect 27196 37508 27252 37564
rect 27252 37508 27256 37564
rect 27192 37504 27256 37508
rect 31952 37564 32016 37568
rect 31952 37508 31956 37564
rect 31956 37508 32012 37564
rect 32012 37508 32016 37564
rect 31952 37504 32016 37508
rect 32032 37564 32096 37568
rect 32032 37508 32036 37564
rect 32036 37508 32092 37564
rect 32092 37508 32096 37564
rect 32032 37504 32096 37508
rect 32112 37564 32176 37568
rect 32112 37508 32116 37564
rect 32116 37508 32172 37564
rect 32172 37508 32176 37564
rect 32112 37504 32176 37508
rect 32192 37564 32256 37568
rect 32192 37508 32196 37564
rect 32196 37508 32252 37564
rect 32252 37508 32256 37564
rect 32192 37504 32256 37508
rect 36952 37564 37016 37568
rect 36952 37508 36956 37564
rect 36956 37508 37012 37564
rect 37012 37508 37016 37564
rect 36952 37504 37016 37508
rect 37032 37564 37096 37568
rect 37032 37508 37036 37564
rect 37036 37508 37092 37564
rect 37092 37508 37096 37564
rect 37032 37504 37096 37508
rect 37112 37564 37176 37568
rect 37112 37508 37116 37564
rect 37116 37508 37172 37564
rect 37172 37508 37176 37564
rect 37112 37504 37176 37508
rect 37192 37564 37256 37568
rect 37192 37508 37196 37564
rect 37196 37508 37252 37564
rect 37252 37508 37256 37564
rect 37192 37504 37256 37508
rect 2612 37020 2676 37024
rect 2612 36964 2616 37020
rect 2616 36964 2672 37020
rect 2672 36964 2676 37020
rect 2612 36960 2676 36964
rect 2692 37020 2756 37024
rect 2692 36964 2696 37020
rect 2696 36964 2752 37020
rect 2752 36964 2756 37020
rect 2692 36960 2756 36964
rect 2772 37020 2836 37024
rect 2772 36964 2776 37020
rect 2776 36964 2832 37020
rect 2832 36964 2836 37020
rect 2772 36960 2836 36964
rect 2852 37020 2916 37024
rect 2852 36964 2856 37020
rect 2856 36964 2912 37020
rect 2912 36964 2916 37020
rect 2852 36960 2916 36964
rect 7612 37020 7676 37024
rect 7612 36964 7616 37020
rect 7616 36964 7672 37020
rect 7672 36964 7676 37020
rect 7612 36960 7676 36964
rect 7692 37020 7756 37024
rect 7692 36964 7696 37020
rect 7696 36964 7752 37020
rect 7752 36964 7756 37020
rect 7692 36960 7756 36964
rect 7772 37020 7836 37024
rect 7772 36964 7776 37020
rect 7776 36964 7832 37020
rect 7832 36964 7836 37020
rect 7772 36960 7836 36964
rect 7852 37020 7916 37024
rect 7852 36964 7856 37020
rect 7856 36964 7912 37020
rect 7912 36964 7916 37020
rect 7852 36960 7916 36964
rect 12612 37020 12676 37024
rect 12612 36964 12616 37020
rect 12616 36964 12672 37020
rect 12672 36964 12676 37020
rect 12612 36960 12676 36964
rect 12692 37020 12756 37024
rect 12692 36964 12696 37020
rect 12696 36964 12752 37020
rect 12752 36964 12756 37020
rect 12692 36960 12756 36964
rect 12772 37020 12836 37024
rect 12772 36964 12776 37020
rect 12776 36964 12832 37020
rect 12832 36964 12836 37020
rect 12772 36960 12836 36964
rect 12852 37020 12916 37024
rect 12852 36964 12856 37020
rect 12856 36964 12912 37020
rect 12912 36964 12916 37020
rect 12852 36960 12916 36964
rect 17612 37020 17676 37024
rect 17612 36964 17616 37020
rect 17616 36964 17672 37020
rect 17672 36964 17676 37020
rect 17612 36960 17676 36964
rect 17692 37020 17756 37024
rect 17692 36964 17696 37020
rect 17696 36964 17752 37020
rect 17752 36964 17756 37020
rect 17692 36960 17756 36964
rect 17772 37020 17836 37024
rect 17772 36964 17776 37020
rect 17776 36964 17832 37020
rect 17832 36964 17836 37020
rect 17772 36960 17836 36964
rect 17852 37020 17916 37024
rect 17852 36964 17856 37020
rect 17856 36964 17912 37020
rect 17912 36964 17916 37020
rect 17852 36960 17916 36964
rect 22612 37020 22676 37024
rect 22612 36964 22616 37020
rect 22616 36964 22672 37020
rect 22672 36964 22676 37020
rect 22612 36960 22676 36964
rect 22692 37020 22756 37024
rect 22692 36964 22696 37020
rect 22696 36964 22752 37020
rect 22752 36964 22756 37020
rect 22692 36960 22756 36964
rect 22772 37020 22836 37024
rect 22772 36964 22776 37020
rect 22776 36964 22832 37020
rect 22832 36964 22836 37020
rect 22772 36960 22836 36964
rect 22852 37020 22916 37024
rect 22852 36964 22856 37020
rect 22856 36964 22912 37020
rect 22912 36964 22916 37020
rect 22852 36960 22916 36964
rect 27612 37020 27676 37024
rect 27612 36964 27616 37020
rect 27616 36964 27672 37020
rect 27672 36964 27676 37020
rect 27612 36960 27676 36964
rect 27692 37020 27756 37024
rect 27692 36964 27696 37020
rect 27696 36964 27752 37020
rect 27752 36964 27756 37020
rect 27692 36960 27756 36964
rect 27772 37020 27836 37024
rect 27772 36964 27776 37020
rect 27776 36964 27832 37020
rect 27832 36964 27836 37020
rect 27772 36960 27836 36964
rect 27852 37020 27916 37024
rect 27852 36964 27856 37020
rect 27856 36964 27912 37020
rect 27912 36964 27916 37020
rect 27852 36960 27916 36964
rect 32612 37020 32676 37024
rect 32612 36964 32616 37020
rect 32616 36964 32672 37020
rect 32672 36964 32676 37020
rect 32612 36960 32676 36964
rect 32692 37020 32756 37024
rect 32692 36964 32696 37020
rect 32696 36964 32752 37020
rect 32752 36964 32756 37020
rect 32692 36960 32756 36964
rect 32772 37020 32836 37024
rect 32772 36964 32776 37020
rect 32776 36964 32832 37020
rect 32832 36964 32836 37020
rect 32772 36960 32836 36964
rect 32852 37020 32916 37024
rect 32852 36964 32856 37020
rect 32856 36964 32912 37020
rect 32912 36964 32916 37020
rect 32852 36960 32916 36964
rect 37612 37020 37676 37024
rect 37612 36964 37616 37020
rect 37616 36964 37672 37020
rect 37672 36964 37676 37020
rect 37612 36960 37676 36964
rect 37692 37020 37756 37024
rect 37692 36964 37696 37020
rect 37696 36964 37752 37020
rect 37752 36964 37756 37020
rect 37692 36960 37756 36964
rect 37772 37020 37836 37024
rect 37772 36964 37776 37020
rect 37776 36964 37832 37020
rect 37832 36964 37836 37020
rect 37772 36960 37836 36964
rect 37852 37020 37916 37024
rect 37852 36964 37856 37020
rect 37856 36964 37912 37020
rect 37912 36964 37916 37020
rect 37852 36960 37916 36964
rect 1952 36476 2016 36480
rect 1952 36420 1956 36476
rect 1956 36420 2012 36476
rect 2012 36420 2016 36476
rect 1952 36416 2016 36420
rect 2032 36476 2096 36480
rect 2032 36420 2036 36476
rect 2036 36420 2092 36476
rect 2092 36420 2096 36476
rect 2032 36416 2096 36420
rect 2112 36476 2176 36480
rect 2112 36420 2116 36476
rect 2116 36420 2172 36476
rect 2172 36420 2176 36476
rect 2112 36416 2176 36420
rect 2192 36476 2256 36480
rect 2192 36420 2196 36476
rect 2196 36420 2252 36476
rect 2252 36420 2256 36476
rect 2192 36416 2256 36420
rect 6952 36476 7016 36480
rect 6952 36420 6956 36476
rect 6956 36420 7012 36476
rect 7012 36420 7016 36476
rect 6952 36416 7016 36420
rect 7032 36476 7096 36480
rect 7032 36420 7036 36476
rect 7036 36420 7092 36476
rect 7092 36420 7096 36476
rect 7032 36416 7096 36420
rect 7112 36476 7176 36480
rect 7112 36420 7116 36476
rect 7116 36420 7172 36476
rect 7172 36420 7176 36476
rect 7112 36416 7176 36420
rect 7192 36476 7256 36480
rect 7192 36420 7196 36476
rect 7196 36420 7252 36476
rect 7252 36420 7256 36476
rect 7192 36416 7256 36420
rect 11952 36476 12016 36480
rect 11952 36420 11956 36476
rect 11956 36420 12012 36476
rect 12012 36420 12016 36476
rect 11952 36416 12016 36420
rect 12032 36476 12096 36480
rect 12032 36420 12036 36476
rect 12036 36420 12092 36476
rect 12092 36420 12096 36476
rect 12032 36416 12096 36420
rect 12112 36476 12176 36480
rect 12112 36420 12116 36476
rect 12116 36420 12172 36476
rect 12172 36420 12176 36476
rect 12112 36416 12176 36420
rect 12192 36476 12256 36480
rect 12192 36420 12196 36476
rect 12196 36420 12252 36476
rect 12252 36420 12256 36476
rect 12192 36416 12256 36420
rect 16952 36476 17016 36480
rect 16952 36420 16956 36476
rect 16956 36420 17012 36476
rect 17012 36420 17016 36476
rect 16952 36416 17016 36420
rect 17032 36476 17096 36480
rect 17032 36420 17036 36476
rect 17036 36420 17092 36476
rect 17092 36420 17096 36476
rect 17032 36416 17096 36420
rect 17112 36476 17176 36480
rect 17112 36420 17116 36476
rect 17116 36420 17172 36476
rect 17172 36420 17176 36476
rect 17112 36416 17176 36420
rect 17192 36476 17256 36480
rect 17192 36420 17196 36476
rect 17196 36420 17252 36476
rect 17252 36420 17256 36476
rect 17192 36416 17256 36420
rect 21952 36476 22016 36480
rect 21952 36420 21956 36476
rect 21956 36420 22012 36476
rect 22012 36420 22016 36476
rect 21952 36416 22016 36420
rect 22032 36476 22096 36480
rect 22032 36420 22036 36476
rect 22036 36420 22092 36476
rect 22092 36420 22096 36476
rect 22032 36416 22096 36420
rect 22112 36476 22176 36480
rect 22112 36420 22116 36476
rect 22116 36420 22172 36476
rect 22172 36420 22176 36476
rect 22112 36416 22176 36420
rect 22192 36476 22256 36480
rect 22192 36420 22196 36476
rect 22196 36420 22252 36476
rect 22252 36420 22256 36476
rect 22192 36416 22256 36420
rect 26952 36476 27016 36480
rect 26952 36420 26956 36476
rect 26956 36420 27012 36476
rect 27012 36420 27016 36476
rect 26952 36416 27016 36420
rect 27032 36476 27096 36480
rect 27032 36420 27036 36476
rect 27036 36420 27092 36476
rect 27092 36420 27096 36476
rect 27032 36416 27096 36420
rect 27112 36476 27176 36480
rect 27112 36420 27116 36476
rect 27116 36420 27172 36476
rect 27172 36420 27176 36476
rect 27112 36416 27176 36420
rect 27192 36476 27256 36480
rect 27192 36420 27196 36476
rect 27196 36420 27252 36476
rect 27252 36420 27256 36476
rect 27192 36416 27256 36420
rect 31952 36476 32016 36480
rect 31952 36420 31956 36476
rect 31956 36420 32012 36476
rect 32012 36420 32016 36476
rect 31952 36416 32016 36420
rect 32032 36476 32096 36480
rect 32032 36420 32036 36476
rect 32036 36420 32092 36476
rect 32092 36420 32096 36476
rect 32032 36416 32096 36420
rect 32112 36476 32176 36480
rect 32112 36420 32116 36476
rect 32116 36420 32172 36476
rect 32172 36420 32176 36476
rect 32112 36416 32176 36420
rect 32192 36476 32256 36480
rect 32192 36420 32196 36476
rect 32196 36420 32252 36476
rect 32252 36420 32256 36476
rect 32192 36416 32256 36420
rect 36952 36476 37016 36480
rect 36952 36420 36956 36476
rect 36956 36420 37012 36476
rect 37012 36420 37016 36476
rect 36952 36416 37016 36420
rect 37032 36476 37096 36480
rect 37032 36420 37036 36476
rect 37036 36420 37092 36476
rect 37092 36420 37096 36476
rect 37032 36416 37096 36420
rect 37112 36476 37176 36480
rect 37112 36420 37116 36476
rect 37116 36420 37172 36476
rect 37172 36420 37176 36476
rect 37112 36416 37176 36420
rect 37192 36476 37256 36480
rect 37192 36420 37196 36476
rect 37196 36420 37252 36476
rect 37252 36420 37256 36476
rect 37192 36416 37256 36420
rect 2612 35932 2676 35936
rect 2612 35876 2616 35932
rect 2616 35876 2672 35932
rect 2672 35876 2676 35932
rect 2612 35872 2676 35876
rect 2692 35932 2756 35936
rect 2692 35876 2696 35932
rect 2696 35876 2752 35932
rect 2752 35876 2756 35932
rect 2692 35872 2756 35876
rect 2772 35932 2836 35936
rect 2772 35876 2776 35932
rect 2776 35876 2832 35932
rect 2832 35876 2836 35932
rect 2772 35872 2836 35876
rect 2852 35932 2916 35936
rect 2852 35876 2856 35932
rect 2856 35876 2912 35932
rect 2912 35876 2916 35932
rect 2852 35872 2916 35876
rect 7612 35932 7676 35936
rect 7612 35876 7616 35932
rect 7616 35876 7672 35932
rect 7672 35876 7676 35932
rect 7612 35872 7676 35876
rect 7692 35932 7756 35936
rect 7692 35876 7696 35932
rect 7696 35876 7752 35932
rect 7752 35876 7756 35932
rect 7692 35872 7756 35876
rect 7772 35932 7836 35936
rect 7772 35876 7776 35932
rect 7776 35876 7832 35932
rect 7832 35876 7836 35932
rect 7772 35872 7836 35876
rect 7852 35932 7916 35936
rect 7852 35876 7856 35932
rect 7856 35876 7912 35932
rect 7912 35876 7916 35932
rect 7852 35872 7916 35876
rect 12612 35932 12676 35936
rect 12612 35876 12616 35932
rect 12616 35876 12672 35932
rect 12672 35876 12676 35932
rect 12612 35872 12676 35876
rect 12692 35932 12756 35936
rect 12692 35876 12696 35932
rect 12696 35876 12752 35932
rect 12752 35876 12756 35932
rect 12692 35872 12756 35876
rect 12772 35932 12836 35936
rect 12772 35876 12776 35932
rect 12776 35876 12832 35932
rect 12832 35876 12836 35932
rect 12772 35872 12836 35876
rect 12852 35932 12916 35936
rect 12852 35876 12856 35932
rect 12856 35876 12912 35932
rect 12912 35876 12916 35932
rect 12852 35872 12916 35876
rect 17612 35932 17676 35936
rect 17612 35876 17616 35932
rect 17616 35876 17672 35932
rect 17672 35876 17676 35932
rect 17612 35872 17676 35876
rect 17692 35932 17756 35936
rect 17692 35876 17696 35932
rect 17696 35876 17752 35932
rect 17752 35876 17756 35932
rect 17692 35872 17756 35876
rect 17772 35932 17836 35936
rect 17772 35876 17776 35932
rect 17776 35876 17832 35932
rect 17832 35876 17836 35932
rect 17772 35872 17836 35876
rect 17852 35932 17916 35936
rect 17852 35876 17856 35932
rect 17856 35876 17912 35932
rect 17912 35876 17916 35932
rect 17852 35872 17916 35876
rect 22612 35932 22676 35936
rect 22612 35876 22616 35932
rect 22616 35876 22672 35932
rect 22672 35876 22676 35932
rect 22612 35872 22676 35876
rect 22692 35932 22756 35936
rect 22692 35876 22696 35932
rect 22696 35876 22752 35932
rect 22752 35876 22756 35932
rect 22692 35872 22756 35876
rect 22772 35932 22836 35936
rect 22772 35876 22776 35932
rect 22776 35876 22832 35932
rect 22832 35876 22836 35932
rect 22772 35872 22836 35876
rect 22852 35932 22916 35936
rect 22852 35876 22856 35932
rect 22856 35876 22912 35932
rect 22912 35876 22916 35932
rect 22852 35872 22916 35876
rect 27612 35932 27676 35936
rect 27612 35876 27616 35932
rect 27616 35876 27672 35932
rect 27672 35876 27676 35932
rect 27612 35872 27676 35876
rect 27692 35932 27756 35936
rect 27692 35876 27696 35932
rect 27696 35876 27752 35932
rect 27752 35876 27756 35932
rect 27692 35872 27756 35876
rect 27772 35932 27836 35936
rect 27772 35876 27776 35932
rect 27776 35876 27832 35932
rect 27832 35876 27836 35932
rect 27772 35872 27836 35876
rect 27852 35932 27916 35936
rect 27852 35876 27856 35932
rect 27856 35876 27912 35932
rect 27912 35876 27916 35932
rect 27852 35872 27916 35876
rect 32612 35932 32676 35936
rect 32612 35876 32616 35932
rect 32616 35876 32672 35932
rect 32672 35876 32676 35932
rect 32612 35872 32676 35876
rect 32692 35932 32756 35936
rect 32692 35876 32696 35932
rect 32696 35876 32752 35932
rect 32752 35876 32756 35932
rect 32692 35872 32756 35876
rect 32772 35932 32836 35936
rect 32772 35876 32776 35932
rect 32776 35876 32832 35932
rect 32832 35876 32836 35932
rect 32772 35872 32836 35876
rect 32852 35932 32916 35936
rect 32852 35876 32856 35932
rect 32856 35876 32912 35932
rect 32912 35876 32916 35932
rect 32852 35872 32916 35876
rect 37612 35932 37676 35936
rect 37612 35876 37616 35932
rect 37616 35876 37672 35932
rect 37672 35876 37676 35932
rect 37612 35872 37676 35876
rect 37692 35932 37756 35936
rect 37692 35876 37696 35932
rect 37696 35876 37752 35932
rect 37752 35876 37756 35932
rect 37692 35872 37756 35876
rect 37772 35932 37836 35936
rect 37772 35876 37776 35932
rect 37776 35876 37832 35932
rect 37832 35876 37836 35932
rect 37772 35872 37836 35876
rect 37852 35932 37916 35936
rect 37852 35876 37856 35932
rect 37856 35876 37912 35932
rect 37912 35876 37916 35932
rect 37852 35872 37916 35876
rect 1952 35388 2016 35392
rect 1952 35332 1956 35388
rect 1956 35332 2012 35388
rect 2012 35332 2016 35388
rect 1952 35328 2016 35332
rect 2032 35388 2096 35392
rect 2032 35332 2036 35388
rect 2036 35332 2092 35388
rect 2092 35332 2096 35388
rect 2032 35328 2096 35332
rect 2112 35388 2176 35392
rect 2112 35332 2116 35388
rect 2116 35332 2172 35388
rect 2172 35332 2176 35388
rect 2112 35328 2176 35332
rect 2192 35388 2256 35392
rect 2192 35332 2196 35388
rect 2196 35332 2252 35388
rect 2252 35332 2256 35388
rect 2192 35328 2256 35332
rect 6952 35388 7016 35392
rect 6952 35332 6956 35388
rect 6956 35332 7012 35388
rect 7012 35332 7016 35388
rect 6952 35328 7016 35332
rect 7032 35388 7096 35392
rect 7032 35332 7036 35388
rect 7036 35332 7092 35388
rect 7092 35332 7096 35388
rect 7032 35328 7096 35332
rect 7112 35388 7176 35392
rect 7112 35332 7116 35388
rect 7116 35332 7172 35388
rect 7172 35332 7176 35388
rect 7112 35328 7176 35332
rect 7192 35388 7256 35392
rect 7192 35332 7196 35388
rect 7196 35332 7252 35388
rect 7252 35332 7256 35388
rect 7192 35328 7256 35332
rect 11952 35388 12016 35392
rect 11952 35332 11956 35388
rect 11956 35332 12012 35388
rect 12012 35332 12016 35388
rect 11952 35328 12016 35332
rect 12032 35388 12096 35392
rect 12032 35332 12036 35388
rect 12036 35332 12092 35388
rect 12092 35332 12096 35388
rect 12032 35328 12096 35332
rect 12112 35388 12176 35392
rect 12112 35332 12116 35388
rect 12116 35332 12172 35388
rect 12172 35332 12176 35388
rect 12112 35328 12176 35332
rect 12192 35388 12256 35392
rect 12192 35332 12196 35388
rect 12196 35332 12252 35388
rect 12252 35332 12256 35388
rect 12192 35328 12256 35332
rect 16952 35388 17016 35392
rect 16952 35332 16956 35388
rect 16956 35332 17012 35388
rect 17012 35332 17016 35388
rect 16952 35328 17016 35332
rect 17032 35388 17096 35392
rect 17032 35332 17036 35388
rect 17036 35332 17092 35388
rect 17092 35332 17096 35388
rect 17032 35328 17096 35332
rect 17112 35388 17176 35392
rect 17112 35332 17116 35388
rect 17116 35332 17172 35388
rect 17172 35332 17176 35388
rect 17112 35328 17176 35332
rect 17192 35388 17256 35392
rect 17192 35332 17196 35388
rect 17196 35332 17252 35388
rect 17252 35332 17256 35388
rect 17192 35328 17256 35332
rect 21952 35388 22016 35392
rect 21952 35332 21956 35388
rect 21956 35332 22012 35388
rect 22012 35332 22016 35388
rect 21952 35328 22016 35332
rect 22032 35388 22096 35392
rect 22032 35332 22036 35388
rect 22036 35332 22092 35388
rect 22092 35332 22096 35388
rect 22032 35328 22096 35332
rect 22112 35388 22176 35392
rect 22112 35332 22116 35388
rect 22116 35332 22172 35388
rect 22172 35332 22176 35388
rect 22112 35328 22176 35332
rect 22192 35388 22256 35392
rect 22192 35332 22196 35388
rect 22196 35332 22252 35388
rect 22252 35332 22256 35388
rect 22192 35328 22256 35332
rect 26952 35388 27016 35392
rect 26952 35332 26956 35388
rect 26956 35332 27012 35388
rect 27012 35332 27016 35388
rect 26952 35328 27016 35332
rect 27032 35388 27096 35392
rect 27032 35332 27036 35388
rect 27036 35332 27092 35388
rect 27092 35332 27096 35388
rect 27032 35328 27096 35332
rect 27112 35388 27176 35392
rect 27112 35332 27116 35388
rect 27116 35332 27172 35388
rect 27172 35332 27176 35388
rect 27112 35328 27176 35332
rect 27192 35388 27256 35392
rect 27192 35332 27196 35388
rect 27196 35332 27252 35388
rect 27252 35332 27256 35388
rect 27192 35328 27256 35332
rect 31952 35388 32016 35392
rect 31952 35332 31956 35388
rect 31956 35332 32012 35388
rect 32012 35332 32016 35388
rect 31952 35328 32016 35332
rect 32032 35388 32096 35392
rect 32032 35332 32036 35388
rect 32036 35332 32092 35388
rect 32092 35332 32096 35388
rect 32032 35328 32096 35332
rect 32112 35388 32176 35392
rect 32112 35332 32116 35388
rect 32116 35332 32172 35388
rect 32172 35332 32176 35388
rect 32112 35328 32176 35332
rect 32192 35388 32256 35392
rect 32192 35332 32196 35388
rect 32196 35332 32252 35388
rect 32252 35332 32256 35388
rect 32192 35328 32256 35332
rect 36952 35388 37016 35392
rect 36952 35332 36956 35388
rect 36956 35332 37012 35388
rect 37012 35332 37016 35388
rect 36952 35328 37016 35332
rect 37032 35388 37096 35392
rect 37032 35332 37036 35388
rect 37036 35332 37092 35388
rect 37092 35332 37096 35388
rect 37032 35328 37096 35332
rect 37112 35388 37176 35392
rect 37112 35332 37116 35388
rect 37116 35332 37172 35388
rect 37172 35332 37176 35388
rect 37112 35328 37176 35332
rect 37192 35388 37256 35392
rect 37192 35332 37196 35388
rect 37196 35332 37252 35388
rect 37252 35332 37256 35388
rect 37192 35328 37256 35332
rect 2612 34844 2676 34848
rect 2612 34788 2616 34844
rect 2616 34788 2672 34844
rect 2672 34788 2676 34844
rect 2612 34784 2676 34788
rect 2692 34844 2756 34848
rect 2692 34788 2696 34844
rect 2696 34788 2752 34844
rect 2752 34788 2756 34844
rect 2692 34784 2756 34788
rect 2772 34844 2836 34848
rect 2772 34788 2776 34844
rect 2776 34788 2832 34844
rect 2832 34788 2836 34844
rect 2772 34784 2836 34788
rect 2852 34844 2916 34848
rect 2852 34788 2856 34844
rect 2856 34788 2912 34844
rect 2912 34788 2916 34844
rect 2852 34784 2916 34788
rect 7612 34844 7676 34848
rect 7612 34788 7616 34844
rect 7616 34788 7672 34844
rect 7672 34788 7676 34844
rect 7612 34784 7676 34788
rect 7692 34844 7756 34848
rect 7692 34788 7696 34844
rect 7696 34788 7752 34844
rect 7752 34788 7756 34844
rect 7692 34784 7756 34788
rect 7772 34844 7836 34848
rect 7772 34788 7776 34844
rect 7776 34788 7832 34844
rect 7832 34788 7836 34844
rect 7772 34784 7836 34788
rect 7852 34844 7916 34848
rect 7852 34788 7856 34844
rect 7856 34788 7912 34844
rect 7912 34788 7916 34844
rect 7852 34784 7916 34788
rect 12612 34844 12676 34848
rect 12612 34788 12616 34844
rect 12616 34788 12672 34844
rect 12672 34788 12676 34844
rect 12612 34784 12676 34788
rect 12692 34844 12756 34848
rect 12692 34788 12696 34844
rect 12696 34788 12752 34844
rect 12752 34788 12756 34844
rect 12692 34784 12756 34788
rect 12772 34844 12836 34848
rect 12772 34788 12776 34844
rect 12776 34788 12832 34844
rect 12832 34788 12836 34844
rect 12772 34784 12836 34788
rect 12852 34844 12916 34848
rect 12852 34788 12856 34844
rect 12856 34788 12912 34844
rect 12912 34788 12916 34844
rect 12852 34784 12916 34788
rect 17612 34844 17676 34848
rect 17612 34788 17616 34844
rect 17616 34788 17672 34844
rect 17672 34788 17676 34844
rect 17612 34784 17676 34788
rect 17692 34844 17756 34848
rect 17692 34788 17696 34844
rect 17696 34788 17752 34844
rect 17752 34788 17756 34844
rect 17692 34784 17756 34788
rect 17772 34844 17836 34848
rect 17772 34788 17776 34844
rect 17776 34788 17832 34844
rect 17832 34788 17836 34844
rect 17772 34784 17836 34788
rect 17852 34844 17916 34848
rect 17852 34788 17856 34844
rect 17856 34788 17912 34844
rect 17912 34788 17916 34844
rect 17852 34784 17916 34788
rect 22612 34844 22676 34848
rect 22612 34788 22616 34844
rect 22616 34788 22672 34844
rect 22672 34788 22676 34844
rect 22612 34784 22676 34788
rect 22692 34844 22756 34848
rect 22692 34788 22696 34844
rect 22696 34788 22752 34844
rect 22752 34788 22756 34844
rect 22692 34784 22756 34788
rect 22772 34844 22836 34848
rect 22772 34788 22776 34844
rect 22776 34788 22832 34844
rect 22832 34788 22836 34844
rect 22772 34784 22836 34788
rect 22852 34844 22916 34848
rect 22852 34788 22856 34844
rect 22856 34788 22912 34844
rect 22912 34788 22916 34844
rect 22852 34784 22916 34788
rect 27612 34844 27676 34848
rect 27612 34788 27616 34844
rect 27616 34788 27672 34844
rect 27672 34788 27676 34844
rect 27612 34784 27676 34788
rect 27692 34844 27756 34848
rect 27692 34788 27696 34844
rect 27696 34788 27752 34844
rect 27752 34788 27756 34844
rect 27692 34784 27756 34788
rect 27772 34844 27836 34848
rect 27772 34788 27776 34844
rect 27776 34788 27832 34844
rect 27832 34788 27836 34844
rect 27772 34784 27836 34788
rect 27852 34844 27916 34848
rect 27852 34788 27856 34844
rect 27856 34788 27912 34844
rect 27912 34788 27916 34844
rect 27852 34784 27916 34788
rect 32612 34844 32676 34848
rect 32612 34788 32616 34844
rect 32616 34788 32672 34844
rect 32672 34788 32676 34844
rect 32612 34784 32676 34788
rect 32692 34844 32756 34848
rect 32692 34788 32696 34844
rect 32696 34788 32752 34844
rect 32752 34788 32756 34844
rect 32692 34784 32756 34788
rect 32772 34844 32836 34848
rect 32772 34788 32776 34844
rect 32776 34788 32832 34844
rect 32832 34788 32836 34844
rect 32772 34784 32836 34788
rect 32852 34844 32916 34848
rect 32852 34788 32856 34844
rect 32856 34788 32912 34844
rect 32912 34788 32916 34844
rect 32852 34784 32916 34788
rect 37612 34844 37676 34848
rect 37612 34788 37616 34844
rect 37616 34788 37672 34844
rect 37672 34788 37676 34844
rect 37612 34784 37676 34788
rect 37692 34844 37756 34848
rect 37692 34788 37696 34844
rect 37696 34788 37752 34844
rect 37752 34788 37756 34844
rect 37692 34784 37756 34788
rect 37772 34844 37836 34848
rect 37772 34788 37776 34844
rect 37776 34788 37832 34844
rect 37832 34788 37836 34844
rect 37772 34784 37836 34788
rect 37852 34844 37916 34848
rect 37852 34788 37856 34844
rect 37856 34788 37912 34844
rect 37912 34788 37916 34844
rect 37852 34784 37916 34788
rect 1952 34300 2016 34304
rect 1952 34244 1956 34300
rect 1956 34244 2012 34300
rect 2012 34244 2016 34300
rect 1952 34240 2016 34244
rect 2032 34300 2096 34304
rect 2032 34244 2036 34300
rect 2036 34244 2092 34300
rect 2092 34244 2096 34300
rect 2032 34240 2096 34244
rect 2112 34300 2176 34304
rect 2112 34244 2116 34300
rect 2116 34244 2172 34300
rect 2172 34244 2176 34300
rect 2112 34240 2176 34244
rect 2192 34300 2256 34304
rect 2192 34244 2196 34300
rect 2196 34244 2252 34300
rect 2252 34244 2256 34300
rect 2192 34240 2256 34244
rect 6952 34300 7016 34304
rect 6952 34244 6956 34300
rect 6956 34244 7012 34300
rect 7012 34244 7016 34300
rect 6952 34240 7016 34244
rect 7032 34300 7096 34304
rect 7032 34244 7036 34300
rect 7036 34244 7092 34300
rect 7092 34244 7096 34300
rect 7032 34240 7096 34244
rect 7112 34300 7176 34304
rect 7112 34244 7116 34300
rect 7116 34244 7172 34300
rect 7172 34244 7176 34300
rect 7112 34240 7176 34244
rect 7192 34300 7256 34304
rect 7192 34244 7196 34300
rect 7196 34244 7252 34300
rect 7252 34244 7256 34300
rect 7192 34240 7256 34244
rect 11952 34300 12016 34304
rect 11952 34244 11956 34300
rect 11956 34244 12012 34300
rect 12012 34244 12016 34300
rect 11952 34240 12016 34244
rect 12032 34300 12096 34304
rect 12032 34244 12036 34300
rect 12036 34244 12092 34300
rect 12092 34244 12096 34300
rect 12032 34240 12096 34244
rect 12112 34300 12176 34304
rect 12112 34244 12116 34300
rect 12116 34244 12172 34300
rect 12172 34244 12176 34300
rect 12112 34240 12176 34244
rect 12192 34300 12256 34304
rect 12192 34244 12196 34300
rect 12196 34244 12252 34300
rect 12252 34244 12256 34300
rect 12192 34240 12256 34244
rect 16952 34300 17016 34304
rect 16952 34244 16956 34300
rect 16956 34244 17012 34300
rect 17012 34244 17016 34300
rect 16952 34240 17016 34244
rect 17032 34300 17096 34304
rect 17032 34244 17036 34300
rect 17036 34244 17092 34300
rect 17092 34244 17096 34300
rect 17032 34240 17096 34244
rect 17112 34300 17176 34304
rect 17112 34244 17116 34300
rect 17116 34244 17172 34300
rect 17172 34244 17176 34300
rect 17112 34240 17176 34244
rect 17192 34300 17256 34304
rect 17192 34244 17196 34300
rect 17196 34244 17252 34300
rect 17252 34244 17256 34300
rect 17192 34240 17256 34244
rect 21952 34300 22016 34304
rect 21952 34244 21956 34300
rect 21956 34244 22012 34300
rect 22012 34244 22016 34300
rect 21952 34240 22016 34244
rect 22032 34300 22096 34304
rect 22032 34244 22036 34300
rect 22036 34244 22092 34300
rect 22092 34244 22096 34300
rect 22032 34240 22096 34244
rect 22112 34300 22176 34304
rect 22112 34244 22116 34300
rect 22116 34244 22172 34300
rect 22172 34244 22176 34300
rect 22112 34240 22176 34244
rect 22192 34300 22256 34304
rect 22192 34244 22196 34300
rect 22196 34244 22252 34300
rect 22252 34244 22256 34300
rect 22192 34240 22256 34244
rect 26952 34300 27016 34304
rect 26952 34244 26956 34300
rect 26956 34244 27012 34300
rect 27012 34244 27016 34300
rect 26952 34240 27016 34244
rect 27032 34300 27096 34304
rect 27032 34244 27036 34300
rect 27036 34244 27092 34300
rect 27092 34244 27096 34300
rect 27032 34240 27096 34244
rect 27112 34300 27176 34304
rect 27112 34244 27116 34300
rect 27116 34244 27172 34300
rect 27172 34244 27176 34300
rect 27112 34240 27176 34244
rect 27192 34300 27256 34304
rect 27192 34244 27196 34300
rect 27196 34244 27252 34300
rect 27252 34244 27256 34300
rect 27192 34240 27256 34244
rect 31952 34300 32016 34304
rect 31952 34244 31956 34300
rect 31956 34244 32012 34300
rect 32012 34244 32016 34300
rect 31952 34240 32016 34244
rect 32032 34300 32096 34304
rect 32032 34244 32036 34300
rect 32036 34244 32092 34300
rect 32092 34244 32096 34300
rect 32032 34240 32096 34244
rect 32112 34300 32176 34304
rect 32112 34244 32116 34300
rect 32116 34244 32172 34300
rect 32172 34244 32176 34300
rect 32112 34240 32176 34244
rect 32192 34300 32256 34304
rect 32192 34244 32196 34300
rect 32196 34244 32252 34300
rect 32252 34244 32256 34300
rect 32192 34240 32256 34244
rect 36952 34300 37016 34304
rect 36952 34244 36956 34300
rect 36956 34244 37012 34300
rect 37012 34244 37016 34300
rect 36952 34240 37016 34244
rect 37032 34300 37096 34304
rect 37032 34244 37036 34300
rect 37036 34244 37092 34300
rect 37092 34244 37096 34300
rect 37032 34240 37096 34244
rect 37112 34300 37176 34304
rect 37112 34244 37116 34300
rect 37116 34244 37172 34300
rect 37172 34244 37176 34300
rect 37112 34240 37176 34244
rect 37192 34300 37256 34304
rect 37192 34244 37196 34300
rect 37196 34244 37252 34300
rect 37252 34244 37256 34300
rect 37192 34240 37256 34244
rect 2612 33756 2676 33760
rect 2612 33700 2616 33756
rect 2616 33700 2672 33756
rect 2672 33700 2676 33756
rect 2612 33696 2676 33700
rect 2692 33756 2756 33760
rect 2692 33700 2696 33756
rect 2696 33700 2752 33756
rect 2752 33700 2756 33756
rect 2692 33696 2756 33700
rect 2772 33756 2836 33760
rect 2772 33700 2776 33756
rect 2776 33700 2832 33756
rect 2832 33700 2836 33756
rect 2772 33696 2836 33700
rect 2852 33756 2916 33760
rect 2852 33700 2856 33756
rect 2856 33700 2912 33756
rect 2912 33700 2916 33756
rect 2852 33696 2916 33700
rect 7612 33756 7676 33760
rect 7612 33700 7616 33756
rect 7616 33700 7672 33756
rect 7672 33700 7676 33756
rect 7612 33696 7676 33700
rect 7692 33756 7756 33760
rect 7692 33700 7696 33756
rect 7696 33700 7752 33756
rect 7752 33700 7756 33756
rect 7692 33696 7756 33700
rect 7772 33756 7836 33760
rect 7772 33700 7776 33756
rect 7776 33700 7832 33756
rect 7832 33700 7836 33756
rect 7772 33696 7836 33700
rect 7852 33756 7916 33760
rect 7852 33700 7856 33756
rect 7856 33700 7912 33756
rect 7912 33700 7916 33756
rect 7852 33696 7916 33700
rect 12612 33756 12676 33760
rect 12612 33700 12616 33756
rect 12616 33700 12672 33756
rect 12672 33700 12676 33756
rect 12612 33696 12676 33700
rect 12692 33756 12756 33760
rect 12692 33700 12696 33756
rect 12696 33700 12752 33756
rect 12752 33700 12756 33756
rect 12692 33696 12756 33700
rect 12772 33756 12836 33760
rect 12772 33700 12776 33756
rect 12776 33700 12832 33756
rect 12832 33700 12836 33756
rect 12772 33696 12836 33700
rect 12852 33756 12916 33760
rect 12852 33700 12856 33756
rect 12856 33700 12912 33756
rect 12912 33700 12916 33756
rect 12852 33696 12916 33700
rect 17612 33756 17676 33760
rect 17612 33700 17616 33756
rect 17616 33700 17672 33756
rect 17672 33700 17676 33756
rect 17612 33696 17676 33700
rect 17692 33756 17756 33760
rect 17692 33700 17696 33756
rect 17696 33700 17752 33756
rect 17752 33700 17756 33756
rect 17692 33696 17756 33700
rect 17772 33756 17836 33760
rect 17772 33700 17776 33756
rect 17776 33700 17832 33756
rect 17832 33700 17836 33756
rect 17772 33696 17836 33700
rect 17852 33756 17916 33760
rect 17852 33700 17856 33756
rect 17856 33700 17912 33756
rect 17912 33700 17916 33756
rect 17852 33696 17916 33700
rect 22612 33756 22676 33760
rect 22612 33700 22616 33756
rect 22616 33700 22672 33756
rect 22672 33700 22676 33756
rect 22612 33696 22676 33700
rect 22692 33756 22756 33760
rect 22692 33700 22696 33756
rect 22696 33700 22752 33756
rect 22752 33700 22756 33756
rect 22692 33696 22756 33700
rect 22772 33756 22836 33760
rect 22772 33700 22776 33756
rect 22776 33700 22832 33756
rect 22832 33700 22836 33756
rect 22772 33696 22836 33700
rect 22852 33756 22916 33760
rect 22852 33700 22856 33756
rect 22856 33700 22912 33756
rect 22912 33700 22916 33756
rect 22852 33696 22916 33700
rect 27612 33756 27676 33760
rect 27612 33700 27616 33756
rect 27616 33700 27672 33756
rect 27672 33700 27676 33756
rect 27612 33696 27676 33700
rect 27692 33756 27756 33760
rect 27692 33700 27696 33756
rect 27696 33700 27752 33756
rect 27752 33700 27756 33756
rect 27692 33696 27756 33700
rect 27772 33756 27836 33760
rect 27772 33700 27776 33756
rect 27776 33700 27832 33756
rect 27832 33700 27836 33756
rect 27772 33696 27836 33700
rect 27852 33756 27916 33760
rect 27852 33700 27856 33756
rect 27856 33700 27912 33756
rect 27912 33700 27916 33756
rect 27852 33696 27916 33700
rect 32612 33756 32676 33760
rect 32612 33700 32616 33756
rect 32616 33700 32672 33756
rect 32672 33700 32676 33756
rect 32612 33696 32676 33700
rect 32692 33756 32756 33760
rect 32692 33700 32696 33756
rect 32696 33700 32752 33756
rect 32752 33700 32756 33756
rect 32692 33696 32756 33700
rect 32772 33756 32836 33760
rect 32772 33700 32776 33756
rect 32776 33700 32832 33756
rect 32832 33700 32836 33756
rect 32772 33696 32836 33700
rect 32852 33756 32916 33760
rect 32852 33700 32856 33756
rect 32856 33700 32912 33756
rect 32912 33700 32916 33756
rect 32852 33696 32916 33700
rect 37612 33756 37676 33760
rect 37612 33700 37616 33756
rect 37616 33700 37672 33756
rect 37672 33700 37676 33756
rect 37612 33696 37676 33700
rect 37692 33756 37756 33760
rect 37692 33700 37696 33756
rect 37696 33700 37752 33756
rect 37752 33700 37756 33756
rect 37692 33696 37756 33700
rect 37772 33756 37836 33760
rect 37772 33700 37776 33756
rect 37776 33700 37832 33756
rect 37832 33700 37836 33756
rect 37772 33696 37836 33700
rect 37852 33756 37916 33760
rect 37852 33700 37856 33756
rect 37856 33700 37912 33756
rect 37912 33700 37916 33756
rect 37852 33696 37916 33700
rect 1952 33212 2016 33216
rect 1952 33156 1956 33212
rect 1956 33156 2012 33212
rect 2012 33156 2016 33212
rect 1952 33152 2016 33156
rect 2032 33212 2096 33216
rect 2032 33156 2036 33212
rect 2036 33156 2092 33212
rect 2092 33156 2096 33212
rect 2032 33152 2096 33156
rect 2112 33212 2176 33216
rect 2112 33156 2116 33212
rect 2116 33156 2172 33212
rect 2172 33156 2176 33212
rect 2112 33152 2176 33156
rect 2192 33212 2256 33216
rect 2192 33156 2196 33212
rect 2196 33156 2252 33212
rect 2252 33156 2256 33212
rect 2192 33152 2256 33156
rect 6952 33212 7016 33216
rect 6952 33156 6956 33212
rect 6956 33156 7012 33212
rect 7012 33156 7016 33212
rect 6952 33152 7016 33156
rect 7032 33212 7096 33216
rect 7032 33156 7036 33212
rect 7036 33156 7092 33212
rect 7092 33156 7096 33212
rect 7032 33152 7096 33156
rect 7112 33212 7176 33216
rect 7112 33156 7116 33212
rect 7116 33156 7172 33212
rect 7172 33156 7176 33212
rect 7112 33152 7176 33156
rect 7192 33212 7256 33216
rect 7192 33156 7196 33212
rect 7196 33156 7252 33212
rect 7252 33156 7256 33212
rect 7192 33152 7256 33156
rect 11952 33212 12016 33216
rect 11952 33156 11956 33212
rect 11956 33156 12012 33212
rect 12012 33156 12016 33212
rect 11952 33152 12016 33156
rect 12032 33212 12096 33216
rect 12032 33156 12036 33212
rect 12036 33156 12092 33212
rect 12092 33156 12096 33212
rect 12032 33152 12096 33156
rect 12112 33212 12176 33216
rect 12112 33156 12116 33212
rect 12116 33156 12172 33212
rect 12172 33156 12176 33212
rect 12112 33152 12176 33156
rect 12192 33212 12256 33216
rect 12192 33156 12196 33212
rect 12196 33156 12252 33212
rect 12252 33156 12256 33212
rect 12192 33152 12256 33156
rect 16952 33212 17016 33216
rect 16952 33156 16956 33212
rect 16956 33156 17012 33212
rect 17012 33156 17016 33212
rect 16952 33152 17016 33156
rect 17032 33212 17096 33216
rect 17032 33156 17036 33212
rect 17036 33156 17092 33212
rect 17092 33156 17096 33212
rect 17032 33152 17096 33156
rect 17112 33212 17176 33216
rect 17112 33156 17116 33212
rect 17116 33156 17172 33212
rect 17172 33156 17176 33212
rect 17112 33152 17176 33156
rect 17192 33212 17256 33216
rect 17192 33156 17196 33212
rect 17196 33156 17252 33212
rect 17252 33156 17256 33212
rect 17192 33152 17256 33156
rect 21952 33212 22016 33216
rect 21952 33156 21956 33212
rect 21956 33156 22012 33212
rect 22012 33156 22016 33212
rect 21952 33152 22016 33156
rect 22032 33212 22096 33216
rect 22032 33156 22036 33212
rect 22036 33156 22092 33212
rect 22092 33156 22096 33212
rect 22032 33152 22096 33156
rect 22112 33212 22176 33216
rect 22112 33156 22116 33212
rect 22116 33156 22172 33212
rect 22172 33156 22176 33212
rect 22112 33152 22176 33156
rect 22192 33212 22256 33216
rect 22192 33156 22196 33212
rect 22196 33156 22252 33212
rect 22252 33156 22256 33212
rect 22192 33152 22256 33156
rect 26952 33212 27016 33216
rect 26952 33156 26956 33212
rect 26956 33156 27012 33212
rect 27012 33156 27016 33212
rect 26952 33152 27016 33156
rect 27032 33212 27096 33216
rect 27032 33156 27036 33212
rect 27036 33156 27092 33212
rect 27092 33156 27096 33212
rect 27032 33152 27096 33156
rect 27112 33212 27176 33216
rect 27112 33156 27116 33212
rect 27116 33156 27172 33212
rect 27172 33156 27176 33212
rect 27112 33152 27176 33156
rect 27192 33212 27256 33216
rect 27192 33156 27196 33212
rect 27196 33156 27252 33212
rect 27252 33156 27256 33212
rect 27192 33152 27256 33156
rect 31952 33212 32016 33216
rect 31952 33156 31956 33212
rect 31956 33156 32012 33212
rect 32012 33156 32016 33212
rect 31952 33152 32016 33156
rect 32032 33212 32096 33216
rect 32032 33156 32036 33212
rect 32036 33156 32092 33212
rect 32092 33156 32096 33212
rect 32032 33152 32096 33156
rect 32112 33212 32176 33216
rect 32112 33156 32116 33212
rect 32116 33156 32172 33212
rect 32172 33156 32176 33212
rect 32112 33152 32176 33156
rect 32192 33212 32256 33216
rect 32192 33156 32196 33212
rect 32196 33156 32252 33212
rect 32252 33156 32256 33212
rect 32192 33152 32256 33156
rect 36952 33212 37016 33216
rect 36952 33156 36956 33212
rect 36956 33156 37012 33212
rect 37012 33156 37016 33212
rect 36952 33152 37016 33156
rect 37032 33212 37096 33216
rect 37032 33156 37036 33212
rect 37036 33156 37092 33212
rect 37092 33156 37096 33212
rect 37032 33152 37096 33156
rect 37112 33212 37176 33216
rect 37112 33156 37116 33212
rect 37116 33156 37172 33212
rect 37172 33156 37176 33212
rect 37112 33152 37176 33156
rect 37192 33212 37256 33216
rect 37192 33156 37196 33212
rect 37196 33156 37252 33212
rect 37252 33156 37256 33212
rect 37192 33152 37256 33156
rect 2612 32668 2676 32672
rect 2612 32612 2616 32668
rect 2616 32612 2672 32668
rect 2672 32612 2676 32668
rect 2612 32608 2676 32612
rect 2692 32668 2756 32672
rect 2692 32612 2696 32668
rect 2696 32612 2752 32668
rect 2752 32612 2756 32668
rect 2692 32608 2756 32612
rect 2772 32668 2836 32672
rect 2772 32612 2776 32668
rect 2776 32612 2832 32668
rect 2832 32612 2836 32668
rect 2772 32608 2836 32612
rect 2852 32668 2916 32672
rect 2852 32612 2856 32668
rect 2856 32612 2912 32668
rect 2912 32612 2916 32668
rect 2852 32608 2916 32612
rect 7612 32668 7676 32672
rect 7612 32612 7616 32668
rect 7616 32612 7672 32668
rect 7672 32612 7676 32668
rect 7612 32608 7676 32612
rect 7692 32668 7756 32672
rect 7692 32612 7696 32668
rect 7696 32612 7752 32668
rect 7752 32612 7756 32668
rect 7692 32608 7756 32612
rect 7772 32668 7836 32672
rect 7772 32612 7776 32668
rect 7776 32612 7832 32668
rect 7832 32612 7836 32668
rect 7772 32608 7836 32612
rect 7852 32668 7916 32672
rect 7852 32612 7856 32668
rect 7856 32612 7912 32668
rect 7912 32612 7916 32668
rect 7852 32608 7916 32612
rect 12612 32668 12676 32672
rect 12612 32612 12616 32668
rect 12616 32612 12672 32668
rect 12672 32612 12676 32668
rect 12612 32608 12676 32612
rect 12692 32668 12756 32672
rect 12692 32612 12696 32668
rect 12696 32612 12752 32668
rect 12752 32612 12756 32668
rect 12692 32608 12756 32612
rect 12772 32668 12836 32672
rect 12772 32612 12776 32668
rect 12776 32612 12832 32668
rect 12832 32612 12836 32668
rect 12772 32608 12836 32612
rect 12852 32668 12916 32672
rect 12852 32612 12856 32668
rect 12856 32612 12912 32668
rect 12912 32612 12916 32668
rect 12852 32608 12916 32612
rect 17612 32668 17676 32672
rect 17612 32612 17616 32668
rect 17616 32612 17672 32668
rect 17672 32612 17676 32668
rect 17612 32608 17676 32612
rect 17692 32668 17756 32672
rect 17692 32612 17696 32668
rect 17696 32612 17752 32668
rect 17752 32612 17756 32668
rect 17692 32608 17756 32612
rect 17772 32668 17836 32672
rect 17772 32612 17776 32668
rect 17776 32612 17832 32668
rect 17832 32612 17836 32668
rect 17772 32608 17836 32612
rect 17852 32668 17916 32672
rect 17852 32612 17856 32668
rect 17856 32612 17912 32668
rect 17912 32612 17916 32668
rect 17852 32608 17916 32612
rect 22612 32668 22676 32672
rect 22612 32612 22616 32668
rect 22616 32612 22672 32668
rect 22672 32612 22676 32668
rect 22612 32608 22676 32612
rect 22692 32668 22756 32672
rect 22692 32612 22696 32668
rect 22696 32612 22752 32668
rect 22752 32612 22756 32668
rect 22692 32608 22756 32612
rect 22772 32668 22836 32672
rect 22772 32612 22776 32668
rect 22776 32612 22832 32668
rect 22832 32612 22836 32668
rect 22772 32608 22836 32612
rect 22852 32668 22916 32672
rect 22852 32612 22856 32668
rect 22856 32612 22912 32668
rect 22912 32612 22916 32668
rect 22852 32608 22916 32612
rect 27612 32668 27676 32672
rect 27612 32612 27616 32668
rect 27616 32612 27672 32668
rect 27672 32612 27676 32668
rect 27612 32608 27676 32612
rect 27692 32668 27756 32672
rect 27692 32612 27696 32668
rect 27696 32612 27752 32668
rect 27752 32612 27756 32668
rect 27692 32608 27756 32612
rect 27772 32668 27836 32672
rect 27772 32612 27776 32668
rect 27776 32612 27832 32668
rect 27832 32612 27836 32668
rect 27772 32608 27836 32612
rect 27852 32668 27916 32672
rect 27852 32612 27856 32668
rect 27856 32612 27912 32668
rect 27912 32612 27916 32668
rect 27852 32608 27916 32612
rect 32612 32668 32676 32672
rect 32612 32612 32616 32668
rect 32616 32612 32672 32668
rect 32672 32612 32676 32668
rect 32612 32608 32676 32612
rect 32692 32668 32756 32672
rect 32692 32612 32696 32668
rect 32696 32612 32752 32668
rect 32752 32612 32756 32668
rect 32692 32608 32756 32612
rect 32772 32668 32836 32672
rect 32772 32612 32776 32668
rect 32776 32612 32832 32668
rect 32832 32612 32836 32668
rect 32772 32608 32836 32612
rect 32852 32668 32916 32672
rect 32852 32612 32856 32668
rect 32856 32612 32912 32668
rect 32912 32612 32916 32668
rect 32852 32608 32916 32612
rect 37612 32668 37676 32672
rect 37612 32612 37616 32668
rect 37616 32612 37672 32668
rect 37672 32612 37676 32668
rect 37612 32608 37676 32612
rect 37692 32668 37756 32672
rect 37692 32612 37696 32668
rect 37696 32612 37752 32668
rect 37752 32612 37756 32668
rect 37692 32608 37756 32612
rect 37772 32668 37836 32672
rect 37772 32612 37776 32668
rect 37776 32612 37832 32668
rect 37832 32612 37836 32668
rect 37772 32608 37836 32612
rect 37852 32668 37916 32672
rect 37852 32612 37856 32668
rect 37856 32612 37912 32668
rect 37912 32612 37916 32668
rect 37852 32608 37916 32612
rect 1952 32124 2016 32128
rect 1952 32068 1956 32124
rect 1956 32068 2012 32124
rect 2012 32068 2016 32124
rect 1952 32064 2016 32068
rect 2032 32124 2096 32128
rect 2032 32068 2036 32124
rect 2036 32068 2092 32124
rect 2092 32068 2096 32124
rect 2032 32064 2096 32068
rect 2112 32124 2176 32128
rect 2112 32068 2116 32124
rect 2116 32068 2172 32124
rect 2172 32068 2176 32124
rect 2112 32064 2176 32068
rect 2192 32124 2256 32128
rect 2192 32068 2196 32124
rect 2196 32068 2252 32124
rect 2252 32068 2256 32124
rect 2192 32064 2256 32068
rect 6952 32124 7016 32128
rect 6952 32068 6956 32124
rect 6956 32068 7012 32124
rect 7012 32068 7016 32124
rect 6952 32064 7016 32068
rect 7032 32124 7096 32128
rect 7032 32068 7036 32124
rect 7036 32068 7092 32124
rect 7092 32068 7096 32124
rect 7032 32064 7096 32068
rect 7112 32124 7176 32128
rect 7112 32068 7116 32124
rect 7116 32068 7172 32124
rect 7172 32068 7176 32124
rect 7112 32064 7176 32068
rect 7192 32124 7256 32128
rect 7192 32068 7196 32124
rect 7196 32068 7252 32124
rect 7252 32068 7256 32124
rect 7192 32064 7256 32068
rect 11952 32124 12016 32128
rect 11952 32068 11956 32124
rect 11956 32068 12012 32124
rect 12012 32068 12016 32124
rect 11952 32064 12016 32068
rect 12032 32124 12096 32128
rect 12032 32068 12036 32124
rect 12036 32068 12092 32124
rect 12092 32068 12096 32124
rect 12032 32064 12096 32068
rect 12112 32124 12176 32128
rect 12112 32068 12116 32124
rect 12116 32068 12172 32124
rect 12172 32068 12176 32124
rect 12112 32064 12176 32068
rect 12192 32124 12256 32128
rect 12192 32068 12196 32124
rect 12196 32068 12252 32124
rect 12252 32068 12256 32124
rect 12192 32064 12256 32068
rect 16952 32124 17016 32128
rect 16952 32068 16956 32124
rect 16956 32068 17012 32124
rect 17012 32068 17016 32124
rect 16952 32064 17016 32068
rect 17032 32124 17096 32128
rect 17032 32068 17036 32124
rect 17036 32068 17092 32124
rect 17092 32068 17096 32124
rect 17032 32064 17096 32068
rect 17112 32124 17176 32128
rect 17112 32068 17116 32124
rect 17116 32068 17172 32124
rect 17172 32068 17176 32124
rect 17112 32064 17176 32068
rect 17192 32124 17256 32128
rect 17192 32068 17196 32124
rect 17196 32068 17252 32124
rect 17252 32068 17256 32124
rect 17192 32064 17256 32068
rect 21952 32124 22016 32128
rect 21952 32068 21956 32124
rect 21956 32068 22012 32124
rect 22012 32068 22016 32124
rect 21952 32064 22016 32068
rect 22032 32124 22096 32128
rect 22032 32068 22036 32124
rect 22036 32068 22092 32124
rect 22092 32068 22096 32124
rect 22032 32064 22096 32068
rect 22112 32124 22176 32128
rect 22112 32068 22116 32124
rect 22116 32068 22172 32124
rect 22172 32068 22176 32124
rect 22112 32064 22176 32068
rect 22192 32124 22256 32128
rect 22192 32068 22196 32124
rect 22196 32068 22252 32124
rect 22252 32068 22256 32124
rect 22192 32064 22256 32068
rect 26952 32124 27016 32128
rect 26952 32068 26956 32124
rect 26956 32068 27012 32124
rect 27012 32068 27016 32124
rect 26952 32064 27016 32068
rect 27032 32124 27096 32128
rect 27032 32068 27036 32124
rect 27036 32068 27092 32124
rect 27092 32068 27096 32124
rect 27032 32064 27096 32068
rect 27112 32124 27176 32128
rect 27112 32068 27116 32124
rect 27116 32068 27172 32124
rect 27172 32068 27176 32124
rect 27112 32064 27176 32068
rect 27192 32124 27256 32128
rect 27192 32068 27196 32124
rect 27196 32068 27252 32124
rect 27252 32068 27256 32124
rect 27192 32064 27256 32068
rect 31952 32124 32016 32128
rect 31952 32068 31956 32124
rect 31956 32068 32012 32124
rect 32012 32068 32016 32124
rect 31952 32064 32016 32068
rect 32032 32124 32096 32128
rect 32032 32068 32036 32124
rect 32036 32068 32092 32124
rect 32092 32068 32096 32124
rect 32032 32064 32096 32068
rect 32112 32124 32176 32128
rect 32112 32068 32116 32124
rect 32116 32068 32172 32124
rect 32172 32068 32176 32124
rect 32112 32064 32176 32068
rect 32192 32124 32256 32128
rect 32192 32068 32196 32124
rect 32196 32068 32252 32124
rect 32252 32068 32256 32124
rect 32192 32064 32256 32068
rect 36952 32124 37016 32128
rect 36952 32068 36956 32124
rect 36956 32068 37012 32124
rect 37012 32068 37016 32124
rect 36952 32064 37016 32068
rect 37032 32124 37096 32128
rect 37032 32068 37036 32124
rect 37036 32068 37092 32124
rect 37092 32068 37096 32124
rect 37032 32064 37096 32068
rect 37112 32124 37176 32128
rect 37112 32068 37116 32124
rect 37116 32068 37172 32124
rect 37172 32068 37176 32124
rect 37112 32064 37176 32068
rect 37192 32124 37256 32128
rect 37192 32068 37196 32124
rect 37196 32068 37252 32124
rect 37252 32068 37256 32124
rect 37192 32064 37256 32068
rect 2612 31580 2676 31584
rect 2612 31524 2616 31580
rect 2616 31524 2672 31580
rect 2672 31524 2676 31580
rect 2612 31520 2676 31524
rect 2692 31580 2756 31584
rect 2692 31524 2696 31580
rect 2696 31524 2752 31580
rect 2752 31524 2756 31580
rect 2692 31520 2756 31524
rect 2772 31580 2836 31584
rect 2772 31524 2776 31580
rect 2776 31524 2832 31580
rect 2832 31524 2836 31580
rect 2772 31520 2836 31524
rect 2852 31580 2916 31584
rect 2852 31524 2856 31580
rect 2856 31524 2912 31580
rect 2912 31524 2916 31580
rect 2852 31520 2916 31524
rect 7612 31580 7676 31584
rect 7612 31524 7616 31580
rect 7616 31524 7672 31580
rect 7672 31524 7676 31580
rect 7612 31520 7676 31524
rect 7692 31580 7756 31584
rect 7692 31524 7696 31580
rect 7696 31524 7752 31580
rect 7752 31524 7756 31580
rect 7692 31520 7756 31524
rect 7772 31580 7836 31584
rect 7772 31524 7776 31580
rect 7776 31524 7832 31580
rect 7832 31524 7836 31580
rect 7772 31520 7836 31524
rect 7852 31580 7916 31584
rect 7852 31524 7856 31580
rect 7856 31524 7912 31580
rect 7912 31524 7916 31580
rect 7852 31520 7916 31524
rect 12612 31580 12676 31584
rect 12612 31524 12616 31580
rect 12616 31524 12672 31580
rect 12672 31524 12676 31580
rect 12612 31520 12676 31524
rect 12692 31580 12756 31584
rect 12692 31524 12696 31580
rect 12696 31524 12752 31580
rect 12752 31524 12756 31580
rect 12692 31520 12756 31524
rect 12772 31580 12836 31584
rect 12772 31524 12776 31580
rect 12776 31524 12832 31580
rect 12832 31524 12836 31580
rect 12772 31520 12836 31524
rect 12852 31580 12916 31584
rect 12852 31524 12856 31580
rect 12856 31524 12912 31580
rect 12912 31524 12916 31580
rect 12852 31520 12916 31524
rect 17612 31580 17676 31584
rect 17612 31524 17616 31580
rect 17616 31524 17672 31580
rect 17672 31524 17676 31580
rect 17612 31520 17676 31524
rect 17692 31580 17756 31584
rect 17692 31524 17696 31580
rect 17696 31524 17752 31580
rect 17752 31524 17756 31580
rect 17692 31520 17756 31524
rect 17772 31580 17836 31584
rect 17772 31524 17776 31580
rect 17776 31524 17832 31580
rect 17832 31524 17836 31580
rect 17772 31520 17836 31524
rect 17852 31580 17916 31584
rect 17852 31524 17856 31580
rect 17856 31524 17912 31580
rect 17912 31524 17916 31580
rect 17852 31520 17916 31524
rect 22612 31580 22676 31584
rect 22612 31524 22616 31580
rect 22616 31524 22672 31580
rect 22672 31524 22676 31580
rect 22612 31520 22676 31524
rect 22692 31580 22756 31584
rect 22692 31524 22696 31580
rect 22696 31524 22752 31580
rect 22752 31524 22756 31580
rect 22692 31520 22756 31524
rect 22772 31580 22836 31584
rect 22772 31524 22776 31580
rect 22776 31524 22832 31580
rect 22832 31524 22836 31580
rect 22772 31520 22836 31524
rect 22852 31580 22916 31584
rect 22852 31524 22856 31580
rect 22856 31524 22912 31580
rect 22912 31524 22916 31580
rect 22852 31520 22916 31524
rect 27612 31580 27676 31584
rect 27612 31524 27616 31580
rect 27616 31524 27672 31580
rect 27672 31524 27676 31580
rect 27612 31520 27676 31524
rect 27692 31580 27756 31584
rect 27692 31524 27696 31580
rect 27696 31524 27752 31580
rect 27752 31524 27756 31580
rect 27692 31520 27756 31524
rect 27772 31580 27836 31584
rect 27772 31524 27776 31580
rect 27776 31524 27832 31580
rect 27832 31524 27836 31580
rect 27772 31520 27836 31524
rect 27852 31580 27916 31584
rect 27852 31524 27856 31580
rect 27856 31524 27912 31580
rect 27912 31524 27916 31580
rect 27852 31520 27916 31524
rect 32612 31580 32676 31584
rect 32612 31524 32616 31580
rect 32616 31524 32672 31580
rect 32672 31524 32676 31580
rect 32612 31520 32676 31524
rect 32692 31580 32756 31584
rect 32692 31524 32696 31580
rect 32696 31524 32752 31580
rect 32752 31524 32756 31580
rect 32692 31520 32756 31524
rect 32772 31580 32836 31584
rect 32772 31524 32776 31580
rect 32776 31524 32832 31580
rect 32832 31524 32836 31580
rect 32772 31520 32836 31524
rect 32852 31580 32916 31584
rect 32852 31524 32856 31580
rect 32856 31524 32912 31580
rect 32912 31524 32916 31580
rect 32852 31520 32916 31524
rect 37612 31580 37676 31584
rect 37612 31524 37616 31580
rect 37616 31524 37672 31580
rect 37672 31524 37676 31580
rect 37612 31520 37676 31524
rect 37692 31580 37756 31584
rect 37692 31524 37696 31580
rect 37696 31524 37752 31580
rect 37752 31524 37756 31580
rect 37692 31520 37756 31524
rect 37772 31580 37836 31584
rect 37772 31524 37776 31580
rect 37776 31524 37832 31580
rect 37832 31524 37836 31580
rect 37772 31520 37836 31524
rect 37852 31580 37916 31584
rect 37852 31524 37856 31580
rect 37856 31524 37912 31580
rect 37912 31524 37916 31580
rect 37852 31520 37916 31524
rect 1952 31036 2016 31040
rect 1952 30980 1956 31036
rect 1956 30980 2012 31036
rect 2012 30980 2016 31036
rect 1952 30976 2016 30980
rect 2032 31036 2096 31040
rect 2032 30980 2036 31036
rect 2036 30980 2092 31036
rect 2092 30980 2096 31036
rect 2032 30976 2096 30980
rect 2112 31036 2176 31040
rect 2112 30980 2116 31036
rect 2116 30980 2172 31036
rect 2172 30980 2176 31036
rect 2112 30976 2176 30980
rect 2192 31036 2256 31040
rect 2192 30980 2196 31036
rect 2196 30980 2252 31036
rect 2252 30980 2256 31036
rect 2192 30976 2256 30980
rect 6952 31036 7016 31040
rect 6952 30980 6956 31036
rect 6956 30980 7012 31036
rect 7012 30980 7016 31036
rect 6952 30976 7016 30980
rect 7032 31036 7096 31040
rect 7032 30980 7036 31036
rect 7036 30980 7092 31036
rect 7092 30980 7096 31036
rect 7032 30976 7096 30980
rect 7112 31036 7176 31040
rect 7112 30980 7116 31036
rect 7116 30980 7172 31036
rect 7172 30980 7176 31036
rect 7112 30976 7176 30980
rect 7192 31036 7256 31040
rect 7192 30980 7196 31036
rect 7196 30980 7252 31036
rect 7252 30980 7256 31036
rect 7192 30976 7256 30980
rect 11952 31036 12016 31040
rect 11952 30980 11956 31036
rect 11956 30980 12012 31036
rect 12012 30980 12016 31036
rect 11952 30976 12016 30980
rect 12032 31036 12096 31040
rect 12032 30980 12036 31036
rect 12036 30980 12092 31036
rect 12092 30980 12096 31036
rect 12032 30976 12096 30980
rect 12112 31036 12176 31040
rect 12112 30980 12116 31036
rect 12116 30980 12172 31036
rect 12172 30980 12176 31036
rect 12112 30976 12176 30980
rect 12192 31036 12256 31040
rect 12192 30980 12196 31036
rect 12196 30980 12252 31036
rect 12252 30980 12256 31036
rect 12192 30976 12256 30980
rect 16952 31036 17016 31040
rect 16952 30980 16956 31036
rect 16956 30980 17012 31036
rect 17012 30980 17016 31036
rect 16952 30976 17016 30980
rect 17032 31036 17096 31040
rect 17032 30980 17036 31036
rect 17036 30980 17092 31036
rect 17092 30980 17096 31036
rect 17032 30976 17096 30980
rect 17112 31036 17176 31040
rect 17112 30980 17116 31036
rect 17116 30980 17172 31036
rect 17172 30980 17176 31036
rect 17112 30976 17176 30980
rect 17192 31036 17256 31040
rect 17192 30980 17196 31036
rect 17196 30980 17252 31036
rect 17252 30980 17256 31036
rect 17192 30976 17256 30980
rect 21952 31036 22016 31040
rect 21952 30980 21956 31036
rect 21956 30980 22012 31036
rect 22012 30980 22016 31036
rect 21952 30976 22016 30980
rect 22032 31036 22096 31040
rect 22032 30980 22036 31036
rect 22036 30980 22092 31036
rect 22092 30980 22096 31036
rect 22032 30976 22096 30980
rect 22112 31036 22176 31040
rect 22112 30980 22116 31036
rect 22116 30980 22172 31036
rect 22172 30980 22176 31036
rect 22112 30976 22176 30980
rect 22192 31036 22256 31040
rect 22192 30980 22196 31036
rect 22196 30980 22252 31036
rect 22252 30980 22256 31036
rect 22192 30976 22256 30980
rect 26952 31036 27016 31040
rect 26952 30980 26956 31036
rect 26956 30980 27012 31036
rect 27012 30980 27016 31036
rect 26952 30976 27016 30980
rect 27032 31036 27096 31040
rect 27032 30980 27036 31036
rect 27036 30980 27092 31036
rect 27092 30980 27096 31036
rect 27032 30976 27096 30980
rect 27112 31036 27176 31040
rect 27112 30980 27116 31036
rect 27116 30980 27172 31036
rect 27172 30980 27176 31036
rect 27112 30976 27176 30980
rect 27192 31036 27256 31040
rect 27192 30980 27196 31036
rect 27196 30980 27252 31036
rect 27252 30980 27256 31036
rect 27192 30976 27256 30980
rect 31952 31036 32016 31040
rect 31952 30980 31956 31036
rect 31956 30980 32012 31036
rect 32012 30980 32016 31036
rect 31952 30976 32016 30980
rect 32032 31036 32096 31040
rect 32032 30980 32036 31036
rect 32036 30980 32092 31036
rect 32092 30980 32096 31036
rect 32032 30976 32096 30980
rect 32112 31036 32176 31040
rect 32112 30980 32116 31036
rect 32116 30980 32172 31036
rect 32172 30980 32176 31036
rect 32112 30976 32176 30980
rect 32192 31036 32256 31040
rect 32192 30980 32196 31036
rect 32196 30980 32252 31036
rect 32252 30980 32256 31036
rect 32192 30976 32256 30980
rect 36952 31036 37016 31040
rect 36952 30980 36956 31036
rect 36956 30980 37012 31036
rect 37012 30980 37016 31036
rect 36952 30976 37016 30980
rect 37032 31036 37096 31040
rect 37032 30980 37036 31036
rect 37036 30980 37092 31036
rect 37092 30980 37096 31036
rect 37032 30976 37096 30980
rect 37112 31036 37176 31040
rect 37112 30980 37116 31036
rect 37116 30980 37172 31036
rect 37172 30980 37176 31036
rect 37112 30976 37176 30980
rect 37192 31036 37256 31040
rect 37192 30980 37196 31036
rect 37196 30980 37252 31036
rect 37252 30980 37256 31036
rect 37192 30976 37256 30980
rect 2612 30492 2676 30496
rect 2612 30436 2616 30492
rect 2616 30436 2672 30492
rect 2672 30436 2676 30492
rect 2612 30432 2676 30436
rect 2692 30492 2756 30496
rect 2692 30436 2696 30492
rect 2696 30436 2752 30492
rect 2752 30436 2756 30492
rect 2692 30432 2756 30436
rect 2772 30492 2836 30496
rect 2772 30436 2776 30492
rect 2776 30436 2832 30492
rect 2832 30436 2836 30492
rect 2772 30432 2836 30436
rect 2852 30492 2916 30496
rect 2852 30436 2856 30492
rect 2856 30436 2912 30492
rect 2912 30436 2916 30492
rect 2852 30432 2916 30436
rect 7612 30492 7676 30496
rect 7612 30436 7616 30492
rect 7616 30436 7672 30492
rect 7672 30436 7676 30492
rect 7612 30432 7676 30436
rect 7692 30492 7756 30496
rect 7692 30436 7696 30492
rect 7696 30436 7752 30492
rect 7752 30436 7756 30492
rect 7692 30432 7756 30436
rect 7772 30492 7836 30496
rect 7772 30436 7776 30492
rect 7776 30436 7832 30492
rect 7832 30436 7836 30492
rect 7772 30432 7836 30436
rect 7852 30492 7916 30496
rect 7852 30436 7856 30492
rect 7856 30436 7912 30492
rect 7912 30436 7916 30492
rect 7852 30432 7916 30436
rect 12612 30492 12676 30496
rect 12612 30436 12616 30492
rect 12616 30436 12672 30492
rect 12672 30436 12676 30492
rect 12612 30432 12676 30436
rect 12692 30492 12756 30496
rect 12692 30436 12696 30492
rect 12696 30436 12752 30492
rect 12752 30436 12756 30492
rect 12692 30432 12756 30436
rect 12772 30492 12836 30496
rect 12772 30436 12776 30492
rect 12776 30436 12832 30492
rect 12832 30436 12836 30492
rect 12772 30432 12836 30436
rect 12852 30492 12916 30496
rect 12852 30436 12856 30492
rect 12856 30436 12912 30492
rect 12912 30436 12916 30492
rect 12852 30432 12916 30436
rect 17612 30492 17676 30496
rect 17612 30436 17616 30492
rect 17616 30436 17672 30492
rect 17672 30436 17676 30492
rect 17612 30432 17676 30436
rect 17692 30492 17756 30496
rect 17692 30436 17696 30492
rect 17696 30436 17752 30492
rect 17752 30436 17756 30492
rect 17692 30432 17756 30436
rect 17772 30492 17836 30496
rect 17772 30436 17776 30492
rect 17776 30436 17832 30492
rect 17832 30436 17836 30492
rect 17772 30432 17836 30436
rect 17852 30492 17916 30496
rect 17852 30436 17856 30492
rect 17856 30436 17912 30492
rect 17912 30436 17916 30492
rect 17852 30432 17916 30436
rect 22612 30492 22676 30496
rect 22612 30436 22616 30492
rect 22616 30436 22672 30492
rect 22672 30436 22676 30492
rect 22612 30432 22676 30436
rect 22692 30492 22756 30496
rect 22692 30436 22696 30492
rect 22696 30436 22752 30492
rect 22752 30436 22756 30492
rect 22692 30432 22756 30436
rect 22772 30492 22836 30496
rect 22772 30436 22776 30492
rect 22776 30436 22832 30492
rect 22832 30436 22836 30492
rect 22772 30432 22836 30436
rect 22852 30492 22916 30496
rect 22852 30436 22856 30492
rect 22856 30436 22912 30492
rect 22912 30436 22916 30492
rect 22852 30432 22916 30436
rect 27612 30492 27676 30496
rect 27612 30436 27616 30492
rect 27616 30436 27672 30492
rect 27672 30436 27676 30492
rect 27612 30432 27676 30436
rect 27692 30492 27756 30496
rect 27692 30436 27696 30492
rect 27696 30436 27752 30492
rect 27752 30436 27756 30492
rect 27692 30432 27756 30436
rect 27772 30492 27836 30496
rect 27772 30436 27776 30492
rect 27776 30436 27832 30492
rect 27832 30436 27836 30492
rect 27772 30432 27836 30436
rect 27852 30492 27916 30496
rect 27852 30436 27856 30492
rect 27856 30436 27912 30492
rect 27912 30436 27916 30492
rect 27852 30432 27916 30436
rect 32612 30492 32676 30496
rect 32612 30436 32616 30492
rect 32616 30436 32672 30492
rect 32672 30436 32676 30492
rect 32612 30432 32676 30436
rect 32692 30492 32756 30496
rect 32692 30436 32696 30492
rect 32696 30436 32752 30492
rect 32752 30436 32756 30492
rect 32692 30432 32756 30436
rect 32772 30492 32836 30496
rect 32772 30436 32776 30492
rect 32776 30436 32832 30492
rect 32832 30436 32836 30492
rect 32772 30432 32836 30436
rect 32852 30492 32916 30496
rect 32852 30436 32856 30492
rect 32856 30436 32912 30492
rect 32912 30436 32916 30492
rect 32852 30432 32916 30436
rect 37612 30492 37676 30496
rect 37612 30436 37616 30492
rect 37616 30436 37672 30492
rect 37672 30436 37676 30492
rect 37612 30432 37676 30436
rect 37692 30492 37756 30496
rect 37692 30436 37696 30492
rect 37696 30436 37752 30492
rect 37752 30436 37756 30492
rect 37692 30432 37756 30436
rect 37772 30492 37836 30496
rect 37772 30436 37776 30492
rect 37776 30436 37832 30492
rect 37832 30436 37836 30492
rect 37772 30432 37836 30436
rect 37852 30492 37916 30496
rect 37852 30436 37856 30492
rect 37856 30436 37912 30492
rect 37912 30436 37916 30492
rect 37852 30432 37916 30436
rect 1952 29948 2016 29952
rect 1952 29892 1956 29948
rect 1956 29892 2012 29948
rect 2012 29892 2016 29948
rect 1952 29888 2016 29892
rect 2032 29948 2096 29952
rect 2032 29892 2036 29948
rect 2036 29892 2092 29948
rect 2092 29892 2096 29948
rect 2032 29888 2096 29892
rect 2112 29948 2176 29952
rect 2112 29892 2116 29948
rect 2116 29892 2172 29948
rect 2172 29892 2176 29948
rect 2112 29888 2176 29892
rect 2192 29948 2256 29952
rect 2192 29892 2196 29948
rect 2196 29892 2252 29948
rect 2252 29892 2256 29948
rect 2192 29888 2256 29892
rect 6952 29948 7016 29952
rect 6952 29892 6956 29948
rect 6956 29892 7012 29948
rect 7012 29892 7016 29948
rect 6952 29888 7016 29892
rect 7032 29948 7096 29952
rect 7032 29892 7036 29948
rect 7036 29892 7092 29948
rect 7092 29892 7096 29948
rect 7032 29888 7096 29892
rect 7112 29948 7176 29952
rect 7112 29892 7116 29948
rect 7116 29892 7172 29948
rect 7172 29892 7176 29948
rect 7112 29888 7176 29892
rect 7192 29948 7256 29952
rect 7192 29892 7196 29948
rect 7196 29892 7252 29948
rect 7252 29892 7256 29948
rect 7192 29888 7256 29892
rect 11952 29948 12016 29952
rect 11952 29892 11956 29948
rect 11956 29892 12012 29948
rect 12012 29892 12016 29948
rect 11952 29888 12016 29892
rect 12032 29948 12096 29952
rect 12032 29892 12036 29948
rect 12036 29892 12092 29948
rect 12092 29892 12096 29948
rect 12032 29888 12096 29892
rect 12112 29948 12176 29952
rect 12112 29892 12116 29948
rect 12116 29892 12172 29948
rect 12172 29892 12176 29948
rect 12112 29888 12176 29892
rect 12192 29948 12256 29952
rect 12192 29892 12196 29948
rect 12196 29892 12252 29948
rect 12252 29892 12256 29948
rect 12192 29888 12256 29892
rect 16952 29948 17016 29952
rect 16952 29892 16956 29948
rect 16956 29892 17012 29948
rect 17012 29892 17016 29948
rect 16952 29888 17016 29892
rect 17032 29948 17096 29952
rect 17032 29892 17036 29948
rect 17036 29892 17092 29948
rect 17092 29892 17096 29948
rect 17032 29888 17096 29892
rect 17112 29948 17176 29952
rect 17112 29892 17116 29948
rect 17116 29892 17172 29948
rect 17172 29892 17176 29948
rect 17112 29888 17176 29892
rect 17192 29948 17256 29952
rect 17192 29892 17196 29948
rect 17196 29892 17252 29948
rect 17252 29892 17256 29948
rect 17192 29888 17256 29892
rect 21952 29948 22016 29952
rect 21952 29892 21956 29948
rect 21956 29892 22012 29948
rect 22012 29892 22016 29948
rect 21952 29888 22016 29892
rect 22032 29948 22096 29952
rect 22032 29892 22036 29948
rect 22036 29892 22092 29948
rect 22092 29892 22096 29948
rect 22032 29888 22096 29892
rect 22112 29948 22176 29952
rect 22112 29892 22116 29948
rect 22116 29892 22172 29948
rect 22172 29892 22176 29948
rect 22112 29888 22176 29892
rect 22192 29948 22256 29952
rect 22192 29892 22196 29948
rect 22196 29892 22252 29948
rect 22252 29892 22256 29948
rect 22192 29888 22256 29892
rect 26952 29948 27016 29952
rect 26952 29892 26956 29948
rect 26956 29892 27012 29948
rect 27012 29892 27016 29948
rect 26952 29888 27016 29892
rect 27032 29948 27096 29952
rect 27032 29892 27036 29948
rect 27036 29892 27092 29948
rect 27092 29892 27096 29948
rect 27032 29888 27096 29892
rect 27112 29948 27176 29952
rect 27112 29892 27116 29948
rect 27116 29892 27172 29948
rect 27172 29892 27176 29948
rect 27112 29888 27176 29892
rect 27192 29948 27256 29952
rect 27192 29892 27196 29948
rect 27196 29892 27252 29948
rect 27252 29892 27256 29948
rect 27192 29888 27256 29892
rect 31952 29948 32016 29952
rect 31952 29892 31956 29948
rect 31956 29892 32012 29948
rect 32012 29892 32016 29948
rect 31952 29888 32016 29892
rect 32032 29948 32096 29952
rect 32032 29892 32036 29948
rect 32036 29892 32092 29948
rect 32092 29892 32096 29948
rect 32032 29888 32096 29892
rect 32112 29948 32176 29952
rect 32112 29892 32116 29948
rect 32116 29892 32172 29948
rect 32172 29892 32176 29948
rect 32112 29888 32176 29892
rect 32192 29948 32256 29952
rect 32192 29892 32196 29948
rect 32196 29892 32252 29948
rect 32252 29892 32256 29948
rect 32192 29888 32256 29892
rect 36952 29948 37016 29952
rect 36952 29892 36956 29948
rect 36956 29892 37012 29948
rect 37012 29892 37016 29948
rect 36952 29888 37016 29892
rect 37032 29948 37096 29952
rect 37032 29892 37036 29948
rect 37036 29892 37092 29948
rect 37092 29892 37096 29948
rect 37032 29888 37096 29892
rect 37112 29948 37176 29952
rect 37112 29892 37116 29948
rect 37116 29892 37172 29948
rect 37172 29892 37176 29948
rect 37112 29888 37176 29892
rect 37192 29948 37256 29952
rect 37192 29892 37196 29948
rect 37196 29892 37252 29948
rect 37252 29892 37256 29948
rect 37192 29888 37256 29892
rect 2612 29404 2676 29408
rect 2612 29348 2616 29404
rect 2616 29348 2672 29404
rect 2672 29348 2676 29404
rect 2612 29344 2676 29348
rect 2692 29404 2756 29408
rect 2692 29348 2696 29404
rect 2696 29348 2752 29404
rect 2752 29348 2756 29404
rect 2692 29344 2756 29348
rect 2772 29404 2836 29408
rect 2772 29348 2776 29404
rect 2776 29348 2832 29404
rect 2832 29348 2836 29404
rect 2772 29344 2836 29348
rect 2852 29404 2916 29408
rect 2852 29348 2856 29404
rect 2856 29348 2912 29404
rect 2912 29348 2916 29404
rect 2852 29344 2916 29348
rect 7612 29404 7676 29408
rect 7612 29348 7616 29404
rect 7616 29348 7672 29404
rect 7672 29348 7676 29404
rect 7612 29344 7676 29348
rect 7692 29404 7756 29408
rect 7692 29348 7696 29404
rect 7696 29348 7752 29404
rect 7752 29348 7756 29404
rect 7692 29344 7756 29348
rect 7772 29404 7836 29408
rect 7772 29348 7776 29404
rect 7776 29348 7832 29404
rect 7832 29348 7836 29404
rect 7772 29344 7836 29348
rect 7852 29404 7916 29408
rect 7852 29348 7856 29404
rect 7856 29348 7912 29404
rect 7912 29348 7916 29404
rect 7852 29344 7916 29348
rect 12612 29404 12676 29408
rect 12612 29348 12616 29404
rect 12616 29348 12672 29404
rect 12672 29348 12676 29404
rect 12612 29344 12676 29348
rect 12692 29404 12756 29408
rect 12692 29348 12696 29404
rect 12696 29348 12752 29404
rect 12752 29348 12756 29404
rect 12692 29344 12756 29348
rect 12772 29404 12836 29408
rect 12772 29348 12776 29404
rect 12776 29348 12832 29404
rect 12832 29348 12836 29404
rect 12772 29344 12836 29348
rect 12852 29404 12916 29408
rect 12852 29348 12856 29404
rect 12856 29348 12912 29404
rect 12912 29348 12916 29404
rect 12852 29344 12916 29348
rect 17612 29404 17676 29408
rect 17612 29348 17616 29404
rect 17616 29348 17672 29404
rect 17672 29348 17676 29404
rect 17612 29344 17676 29348
rect 17692 29404 17756 29408
rect 17692 29348 17696 29404
rect 17696 29348 17752 29404
rect 17752 29348 17756 29404
rect 17692 29344 17756 29348
rect 17772 29404 17836 29408
rect 17772 29348 17776 29404
rect 17776 29348 17832 29404
rect 17832 29348 17836 29404
rect 17772 29344 17836 29348
rect 17852 29404 17916 29408
rect 17852 29348 17856 29404
rect 17856 29348 17912 29404
rect 17912 29348 17916 29404
rect 17852 29344 17916 29348
rect 22612 29404 22676 29408
rect 22612 29348 22616 29404
rect 22616 29348 22672 29404
rect 22672 29348 22676 29404
rect 22612 29344 22676 29348
rect 22692 29404 22756 29408
rect 22692 29348 22696 29404
rect 22696 29348 22752 29404
rect 22752 29348 22756 29404
rect 22692 29344 22756 29348
rect 22772 29404 22836 29408
rect 22772 29348 22776 29404
rect 22776 29348 22832 29404
rect 22832 29348 22836 29404
rect 22772 29344 22836 29348
rect 22852 29404 22916 29408
rect 22852 29348 22856 29404
rect 22856 29348 22912 29404
rect 22912 29348 22916 29404
rect 22852 29344 22916 29348
rect 27612 29404 27676 29408
rect 27612 29348 27616 29404
rect 27616 29348 27672 29404
rect 27672 29348 27676 29404
rect 27612 29344 27676 29348
rect 27692 29404 27756 29408
rect 27692 29348 27696 29404
rect 27696 29348 27752 29404
rect 27752 29348 27756 29404
rect 27692 29344 27756 29348
rect 27772 29404 27836 29408
rect 27772 29348 27776 29404
rect 27776 29348 27832 29404
rect 27832 29348 27836 29404
rect 27772 29344 27836 29348
rect 27852 29404 27916 29408
rect 27852 29348 27856 29404
rect 27856 29348 27912 29404
rect 27912 29348 27916 29404
rect 27852 29344 27916 29348
rect 32612 29404 32676 29408
rect 32612 29348 32616 29404
rect 32616 29348 32672 29404
rect 32672 29348 32676 29404
rect 32612 29344 32676 29348
rect 32692 29404 32756 29408
rect 32692 29348 32696 29404
rect 32696 29348 32752 29404
rect 32752 29348 32756 29404
rect 32692 29344 32756 29348
rect 32772 29404 32836 29408
rect 32772 29348 32776 29404
rect 32776 29348 32832 29404
rect 32832 29348 32836 29404
rect 32772 29344 32836 29348
rect 32852 29404 32916 29408
rect 32852 29348 32856 29404
rect 32856 29348 32912 29404
rect 32912 29348 32916 29404
rect 32852 29344 32916 29348
rect 37612 29404 37676 29408
rect 37612 29348 37616 29404
rect 37616 29348 37672 29404
rect 37672 29348 37676 29404
rect 37612 29344 37676 29348
rect 37692 29404 37756 29408
rect 37692 29348 37696 29404
rect 37696 29348 37752 29404
rect 37752 29348 37756 29404
rect 37692 29344 37756 29348
rect 37772 29404 37836 29408
rect 37772 29348 37776 29404
rect 37776 29348 37832 29404
rect 37832 29348 37836 29404
rect 37772 29344 37836 29348
rect 37852 29404 37916 29408
rect 37852 29348 37856 29404
rect 37856 29348 37912 29404
rect 37912 29348 37916 29404
rect 37852 29344 37916 29348
rect 1952 28860 2016 28864
rect 1952 28804 1956 28860
rect 1956 28804 2012 28860
rect 2012 28804 2016 28860
rect 1952 28800 2016 28804
rect 2032 28860 2096 28864
rect 2032 28804 2036 28860
rect 2036 28804 2092 28860
rect 2092 28804 2096 28860
rect 2032 28800 2096 28804
rect 2112 28860 2176 28864
rect 2112 28804 2116 28860
rect 2116 28804 2172 28860
rect 2172 28804 2176 28860
rect 2112 28800 2176 28804
rect 2192 28860 2256 28864
rect 2192 28804 2196 28860
rect 2196 28804 2252 28860
rect 2252 28804 2256 28860
rect 2192 28800 2256 28804
rect 6952 28860 7016 28864
rect 6952 28804 6956 28860
rect 6956 28804 7012 28860
rect 7012 28804 7016 28860
rect 6952 28800 7016 28804
rect 7032 28860 7096 28864
rect 7032 28804 7036 28860
rect 7036 28804 7092 28860
rect 7092 28804 7096 28860
rect 7032 28800 7096 28804
rect 7112 28860 7176 28864
rect 7112 28804 7116 28860
rect 7116 28804 7172 28860
rect 7172 28804 7176 28860
rect 7112 28800 7176 28804
rect 7192 28860 7256 28864
rect 7192 28804 7196 28860
rect 7196 28804 7252 28860
rect 7252 28804 7256 28860
rect 7192 28800 7256 28804
rect 11952 28860 12016 28864
rect 11952 28804 11956 28860
rect 11956 28804 12012 28860
rect 12012 28804 12016 28860
rect 11952 28800 12016 28804
rect 12032 28860 12096 28864
rect 12032 28804 12036 28860
rect 12036 28804 12092 28860
rect 12092 28804 12096 28860
rect 12032 28800 12096 28804
rect 12112 28860 12176 28864
rect 12112 28804 12116 28860
rect 12116 28804 12172 28860
rect 12172 28804 12176 28860
rect 12112 28800 12176 28804
rect 12192 28860 12256 28864
rect 12192 28804 12196 28860
rect 12196 28804 12252 28860
rect 12252 28804 12256 28860
rect 12192 28800 12256 28804
rect 16952 28860 17016 28864
rect 16952 28804 16956 28860
rect 16956 28804 17012 28860
rect 17012 28804 17016 28860
rect 16952 28800 17016 28804
rect 17032 28860 17096 28864
rect 17032 28804 17036 28860
rect 17036 28804 17092 28860
rect 17092 28804 17096 28860
rect 17032 28800 17096 28804
rect 17112 28860 17176 28864
rect 17112 28804 17116 28860
rect 17116 28804 17172 28860
rect 17172 28804 17176 28860
rect 17112 28800 17176 28804
rect 17192 28860 17256 28864
rect 17192 28804 17196 28860
rect 17196 28804 17252 28860
rect 17252 28804 17256 28860
rect 17192 28800 17256 28804
rect 21952 28860 22016 28864
rect 21952 28804 21956 28860
rect 21956 28804 22012 28860
rect 22012 28804 22016 28860
rect 21952 28800 22016 28804
rect 22032 28860 22096 28864
rect 22032 28804 22036 28860
rect 22036 28804 22092 28860
rect 22092 28804 22096 28860
rect 22032 28800 22096 28804
rect 22112 28860 22176 28864
rect 22112 28804 22116 28860
rect 22116 28804 22172 28860
rect 22172 28804 22176 28860
rect 22112 28800 22176 28804
rect 22192 28860 22256 28864
rect 22192 28804 22196 28860
rect 22196 28804 22252 28860
rect 22252 28804 22256 28860
rect 22192 28800 22256 28804
rect 26952 28860 27016 28864
rect 26952 28804 26956 28860
rect 26956 28804 27012 28860
rect 27012 28804 27016 28860
rect 26952 28800 27016 28804
rect 27032 28860 27096 28864
rect 27032 28804 27036 28860
rect 27036 28804 27092 28860
rect 27092 28804 27096 28860
rect 27032 28800 27096 28804
rect 27112 28860 27176 28864
rect 27112 28804 27116 28860
rect 27116 28804 27172 28860
rect 27172 28804 27176 28860
rect 27112 28800 27176 28804
rect 27192 28860 27256 28864
rect 27192 28804 27196 28860
rect 27196 28804 27252 28860
rect 27252 28804 27256 28860
rect 27192 28800 27256 28804
rect 31952 28860 32016 28864
rect 31952 28804 31956 28860
rect 31956 28804 32012 28860
rect 32012 28804 32016 28860
rect 31952 28800 32016 28804
rect 32032 28860 32096 28864
rect 32032 28804 32036 28860
rect 32036 28804 32092 28860
rect 32092 28804 32096 28860
rect 32032 28800 32096 28804
rect 32112 28860 32176 28864
rect 32112 28804 32116 28860
rect 32116 28804 32172 28860
rect 32172 28804 32176 28860
rect 32112 28800 32176 28804
rect 32192 28860 32256 28864
rect 32192 28804 32196 28860
rect 32196 28804 32252 28860
rect 32252 28804 32256 28860
rect 32192 28800 32256 28804
rect 36952 28860 37016 28864
rect 36952 28804 36956 28860
rect 36956 28804 37012 28860
rect 37012 28804 37016 28860
rect 36952 28800 37016 28804
rect 37032 28860 37096 28864
rect 37032 28804 37036 28860
rect 37036 28804 37092 28860
rect 37092 28804 37096 28860
rect 37032 28800 37096 28804
rect 37112 28860 37176 28864
rect 37112 28804 37116 28860
rect 37116 28804 37172 28860
rect 37172 28804 37176 28860
rect 37112 28800 37176 28804
rect 37192 28860 37256 28864
rect 37192 28804 37196 28860
rect 37196 28804 37252 28860
rect 37252 28804 37256 28860
rect 37192 28800 37256 28804
rect 2612 28316 2676 28320
rect 2612 28260 2616 28316
rect 2616 28260 2672 28316
rect 2672 28260 2676 28316
rect 2612 28256 2676 28260
rect 2692 28316 2756 28320
rect 2692 28260 2696 28316
rect 2696 28260 2752 28316
rect 2752 28260 2756 28316
rect 2692 28256 2756 28260
rect 2772 28316 2836 28320
rect 2772 28260 2776 28316
rect 2776 28260 2832 28316
rect 2832 28260 2836 28316
rect 2772 28256 2836 28260
rect 2852 28316 2916 28320
rect 2852 28260 2856 28316
rect 2856 28260 2912 28316
rect 2912 28260 2916 28316
rect 2852 28256 2916 28260
rect 7612 28316 7676 28320
rect 7612 28260 7616 28316
rect 7616 28260 7672 28316
rect 7672 28260 7676 28316
rect 7612 28256 7676 28260
rect 7692 28316 7756 28320
rect 7692 28260 7696 28316
rect 7696 28260 7752 28316
rect 7752 28260 7756 28316
rect 7692 28256 7756 28260
rect 7772 28316 7836 28320
rect 7772 28260 7776 28316
rect 7776 28260 7832 28316
rect 7832 28260 7836 28316
rect 7772 28256 7836 28260
rect 7852 28316 7916 28320
rect 7852 28260 7856 28316
rect 7856 28260 7912 28316
rect 7912 28260 7916 28316
rect 7852 28256 7916 28260
rect 12612 28316 12676 28320
rect 12612 28260 12616 28316
rect 12616 28260 12672 28316
rect 12672 28260 12676 28316
rect 12612 28256 12676 28260
rect 12692 28316 12756 28320
rect 12692 28260 12696 28316
rect 12696 28260 12752 28316
rect 12752 28260 12756 28316
rect 12692 28256 12756 28260
rect 12772 28316 12836 28320
rect 12772 28260 12776 28316
rect 12776 28260 12832 28316
rect 12832 28260 12836 28316
rect 12772 28256 12836 28260
rect 12852 28316 12916 28320
rect 12852 28260 12856 28316
rect 12856 28260 12912 28316
rect 12912 28260 12916 28316
rect 12852 28256 12916 28260
rect 17612 28316 17676 28320
rect 17612 28260 17616 28316
rect 17616 28260 17672 28316
rect 17672 28260 17676 28316
rect 17612 28256 17676 28260
rect 17692 28316 17756 28320
rect 17692 28260 17696 28316
rect 17696 28260 17752 28316
rect 17752 28260 17756 28316
rect 17692 28256 17756 28260
rect 17772 28316 17836 28320
rect 17772 28260 17776 28316
rect 17776 28260 17832 28316
rect 17832 28260 17836 28316
rect 17772 28256 17836 28260
rect 17852 28316 17916 28320
rect 17852 28260 17856 28316
rect 17856 28260 17912 28316
rect 17912 28260 17916 28316
rect 17852 28256 17916 28260
rect 22612 28316 22676 28320
rect 22612 28260 22616 28316
rect 22616 28260 22672 28316
rect 22672 28260 22676 28316
rect 22612 28256 22676 28260
rect 22692 28316 22756 28320
rect 22692 28260 22696 28316
rect 22696 28260 22752 28316
rect 22752 28260 22756 28316
rect 22692 28256 22756 28260
rect 22772 28316 22836 28320
rect 22772 28260 22776 28316
rect 22776 28260 22832 28316
rect 22832 28260 22836 28316
rect 22772 28256 22836 28260
rect 22852 28316 22916 28320
rect 22852 28260 22856 28316
rect 22856 28260 22912 28316
rect 22912 28260 22916 28316
rect 22852 28256 22916 28260
rect 27612 28316 27676 28320
rect 27612 28260 27616 28316
rect 27616 28260 27672 28316
rect 27672 28260 27676 28316
rect 27612 28256 27676 28260
rect 27692 28316 27756 28320
rect 27692 28260 27696 28316
rect 27696 28260 27752 28316
rect 27752 28260 27756 28316
rect 27692 28256 27756 28260
rect 27772 28316 27836 28320
rect 27772 28260 27776 28316
rect 27776 28260 27832 28316
rect 27832 28260 27836 28316
rect 27772 28256 27836 28260
rect 27852 28316 27916 28320
rect 27852 28260 27856 28316
rect 27856 28260 27912 28316
rect 27912 28260 27916 28316
rect 27852 28256 27916 28260
rect 32612 28316 32676 28320
rect 32612 28260 32616 28316
rect 32616 28260 32672 28316
rect 32672 28260 32676 28316
rect 32612 28256 32676 28260
rect 32692 28316 32756 28320
rect 32692 28260 32696 28316
rect 32696 28260 32752 28316
rect 32752 28260 32756 28316
rect 32692 28256 32756 28260
rect 32772 28316 32836 28320
rect 32772 28260 32776 28316
rect 32776 28260 32832 28316
rect 32832 28260 32836 28316
rect 32772 28256 32836 28260
rect 32852 28316 32916 28320
rect 32852 28260 32856 28316
rect 32856 28260 32912 28316
rect 32912 28260 32916 28316
rect 32852 28256 32916 28260
rect 37612 28316 37676 28320
rect 37612 28260 37616 28316
rect 37616 28260 37672 28316
rect 37672 28260 37676 28316
rect 37612 28256 37676 28260
rect 37692 28316 37756 28320
rect 37692 28260 37696 28316
rect 37696 28260 37752 28316
rect 37752 28260 37756 28316
rect 37692 28256 37756 28260
rect 37772 28316 37836 28320
rect 37772 28260 37776 28316
rect 37776 28260 37832 28316
rect 37832 28260 37836 28316
rect 37772 28256 37836 28260
rect 37852 28316 37916 28320
rect 37852 28260 37856 28316
rect 37856 28260 37912 28316
rect 37912 28260 37916 28316
rect 37852 28256 37916 28260
rect 1952 27772 2016 27776
rect 1952 27716 1956 27772
rect 1956 27716 2012 27772
rect 2012 27716 2016 27772
rect 1952 27712 2016 27716
rect 2032 27772 2096 27776
rect 2032 27716 2036 27772
rect 2036 27716 2092 27772
rect 2092 27716 2096 27772
rect 2032 27712 2096 27716
rect 2112 27772 2176 27776
rect 2112 27716 2116 27772
rect 2116 27716 2172 27772
rect 2172 27716 2176 27772
rect 2112 27712 2176 27716
rect 2192 27772 2256 27776
rect 2192 27716 2196 27772
rect 2196 27716 2252 27772
rect 2252 27716 2256 27772
rect 2192 27712 2256 27716
rect 6952 27772 7016 27776
rect 6952 27716 6956 27772
rect 6956 27716 7012 27772
rect 7012 27716 7016 27772
rect 6952 27712 7016 27716
rect 7032 27772 7096 27776
rect 7032 27716 7036 27772
rect 7036 27716 7092 27772
rect 7092 27716 7096 27772
rect 7032 27712 7096 27716
rect 7112 27772 7176 27776
rect 7112 27716 7116 27772
rect 7116 27716 7172 27772
rect 7172 27716 7176 27772
rect 7112 27712 7176 27716
rect 7192 27772 7256 27776
rect 7192 27716 7196 27772
rect 7196 27716 7252 27772
rect 7252 27716 7256 27772
rect 7192 27712 7256 27716
rect 11952 27772 12016 27776
rect 11952 27716 11956 27772
rect 11956 27716 12012 27772
rect 12012 27716 12016 27772
rect 11952 27712 12016 27716
rect 12032 27772 12096 27776
rect 12032 27716 12036 27772
rect 12036 27716 12092 27772
rect 12092 27716 12096 27772
rect 12032 27712 12096 27716
rect 12112 27772 12176 27776
rect 12112 27716 12116 27772
rect 12116 27716 12172 27772
rect 12172 27716 12176 27772
rect 12112 27712 12176 27716
rect 12192 27772 12256 27776
rect 12192 27716 12196 27772
rect 12196 27716 12252 27772
rect 12252 27716 12256 27772
rect 12192 27712 12256 27716
rect 16952 27772 17016 27776
rect 16952 27716 16956 27772
rect 16956 27716 17012 27772
rect 17012 27716 17016 27772
rect 16952 27712 17016 27716
rect 17032 27772 17096 27776
rect 17032 27716 17036 27772
rect 17036 27716 17092 27772
rect 17092 27716 17096 27772
rect 17032 27712 17096 27716
rect 17112 27772 17176 27776
rect 17112 27716 17116 27772
rect 17116 27716 17172 27772
rect 17172 27716 17176 27772
rect 17112 27712 17176 27716
rect 17192 27772 17256 27776
rect 17192 27716 17196 27772
rect 17196 27716 17252 27772
rect 17252 27716 17256 27772
rect 17192 27712 17256 27716
rect 21952 27772 22016 27776
rect 21952 27716 21956 27772
rect 21956 27716 22012 27772
rect 22012 27716 22016 27772
rect 21952 27712 22016 27716
rect 22032 27772 22096 27776
rect 22032 27716 22036 27772
rect 22036 27716 22092 27772
rect 22092 27716 22096 27772
rect 22032 27712 22096 27716
rect 22112 27772 22176 27776
rect 22112 27716 22116 27772
rect 22116 27716 22172 27772
rect 22172 27716 22176 27772
rect 22112 27712 22176 27716
rect 22192 27772 22256 27776
rect 22192 27716 22196 27772
rect 22196 27716 22252 27772
rect 22252 27716 22256 27772
rect 22192 27712 22256 27716
rect 26952 27772 27016 27776
rect 26952 27716 26956 27772
rect 26956 27716 27012 27772
rect 27012 27716 27016 27772
rect 26952 27712 27016 27716
rect 27032 27772 27096 27776
rect 27032 27716 27036 27772
rect 27036 27716 27092 27772
rect 27092 27716 27096 27772
rect 27032 27712 27096 27716
rect 27112 27772 27176 27776
rect 27112 27716 27116 27772
rect 27116 27716 27172 27772
rect 27172 27716 27176 27772
rect 27112 27712 27176 27716
rect 27192 27772 27256 27776
rect 27192 27716 27196 27772
rect 27196 27716 27252 27772
rect 27252 27716 27256 27772
rect 27192 27712 27256 27716
rect 31952 27772 32016 27776
rect 31952 27716 31956 27772
rect 31956 27716 32012 27772
rect 32012 27716 32016 27772
rect 31952 27712 32016 27716
rect 32032 27772 32096 27776
rect 32032 27716 32036 27772
rect 32036 27716 32092 27772
rect 32092 27716 32096 27772
rect 32032 27712 32096 27716
rect 32112 27772 32176 27776
rect 32112 27716 32116 27772
rect 32116 27716 32172 27772
rect 32172 27716 32176 27772
rect 32112 27712 32176 27716
rect 32192 27772 32256 27776
rect 32192 27716 32196 27772
rect 32196 27716 32252 27772
rect 32252 27716 32256 27772
rect 32192 27712 32256 27716
rect 36952 27772 37016 27776
rect 36952 27716 36956 27772
rect 36956 27716 37012 27772
rect 37012 27716 37016 27772
rect 36952 27712 37016 27716
rect 37032 27772 37096 27776
rect 37032 27716 37036 27772
rect 37036 27716 37092 27772
rect 37092 27716 37096 27772
rect 37032 27712 37096 27716
rect 37112 27772 37176 27776
rect 37112 27716 37116 27772
rect 37116 27716 37172 27772
rect 37172 27716 37176 27772
rect 37112 27712 37176 27716
rect 37192 27772 37256 27776
rect 37192 27716 37196 27772
rect 37196 27716 37252 27772
rect 37252 27716 37256 27772
rect 37192 27712 37256 27716
rect 2612 27228 2676 27232
rect 2612 27172 2616 27228
rect 2616 27172 2672 27228
rect 2672 27172 2676 27228
rect 2612 27168 2676 27172
rect 2692 27228 2756 27232
rect 2692 27172 2696 27228
rect 2696 27172 2752 27228
rect 2752 27172 2756 27228
rect 2692 27168 2756 27172
rect 2772 27228 2836 27232
rect 2772 27172 2776 27228
rect 2776 27172 2832 27228
rect 2832 27172 2836 27228
rect 2772 27168 2836 27172
rect 2852 27228 2916 27232
rect 2852 27172 2856 27228
rect 2856 27172 2912 27228
rect 2912 27172 2916 27228
rect 2852 27168 2916 27172
rect 7612 27228 7676 27232
rect 7612 27172 7616 27228
rect 7616 27172 7672 27228
rect 7672 27172 7676 27228
rect 7612 27168 7676 27172
rect 7692 27228 7756 27232
rect 7692 27172 7696 27228
rect 7696 27172 7752 27228
rect 7752 27172 7756 27228
rect 7692 27168 7756 27172
rect 7772 27228 7836 27232
rect 7772 27172 7776 27228
rect 7776 27172 7832 27228
rect 7832 27172 7836 27228
rect 7772 27168 7836 27172
rect 7852 27228 7916 27232
rect 7852 27172 7856 27228
rect 7856 27172 7912 27228
rect 7912 27172 7916 27228
rect 7852 27168 7916 27172
rect 12612 27228 12676 27232
rect 12612 27172 12616 27228
rect 12616 27172 12672 27228
rect 12672 27172 12676 27228
rect 12612 27168 12676 27172
rect 12692 27228 12756 27232
rect 12692 27172 12696 27228
rect 12696 27172 12752 27228
rect 12752 27172 12756 27228
rect 12692 27168 12756 27172
rect 12772 27228 12836 27232
rect 12772 27172 12776 27228
rect 12776 27172 12832 27228
rect 12832 27172 12836 27228
rect 12772 27168 12836 27172
rect 12852 27228 12916 27232
rect 12852 27172 12856 27228
rect 12856 27172 12912 27228
rect 12912 27172 12916 27228
rect 12852 27168 12916 27172
rect 17612 27228 17676 27232
rect 17612 27172 17616 27228
rect 17616 27172 17672 27228
rect 17672 27172 17676 27228
rect 17612 27168 17676 27172
rect 17692 27228 17756 27232
rect 17692 27172 17696 27228
rect 17696 27172 17752 27228
rect 17752 27172 17756 27228
rect 17692 27168 17756 27172
rect 17772 27228 17836 27232
rect 17772 27172 17776 27228
rect 17776 27172 17832 27228
rect 17832 27172 17836 27228
rect 17772 27168 17836 27172
rect 17852 27228 17916 27232
rect 17852 27172 17856 27228
rect 17856 27172 17912 27228
rect 17912 27172 17916 27228
rect 17852 27168 17916 27172
rect 22612 27228 22676 27232
rect 22612 27172 22616 27228
rect 22616 27172 22672 27228
rect 22672 27172 22676 27228
rect 22612 27168 22676 27172
rect 22692 27228 22756 27232
rect 22692 27172 22696 27228
rect 22696 27172 22752 27228
rect 22752 27172 22756 27228
rect 22692 27168 22756 27172
rect 22772 27228 22836 27232
rect 22772 27172 22776 27228
rect 22776 27172 22832 27228
rect 22832 27172 22836 27228
rect 22772 27168 22836 27172
rect 22852 27228 22916 27232
rect 22852 27172 22856 27228
rect 22856 27172 22912 27228
rect 22912 27172 22916 27228
rect 22852 27168 22916 27172
rect 27612 27228 27676 27232
rect 27612 27172 27616 27228
rect 27616 27172 27672 27228
rect 27672 27172 27676 27228
rect 27612 27168 27676 27172
rect 27692 27228 27756 27232
rect 27692 27172 27696 27228
rect 27696 27172 27752 27228
rect 27752 27172 27756 27228
rect 27692 27168 27756 27172
rect 27772 27228 27836 27232
rect 27772 27172 27776 27228
rect 27776 27172 27832 27228
rect 27832 27172 27836 27228
rect 27772 27168 27836 27172
rect 27852 27228 27916 27232
rect 27852 27172 27856 27228
rect 27856 27172 27912 27228
rect 27912 27172 27916 27228
rect 27852 27168 27916 27172
rect 32612 27228 32676 27232
rect 32612 27172 32616 27228
rect 32616 27172 32672 27228
rect 32672 27172 32676 27228
rect 32612 27168 32676 27172
rect 32692 27228 32756 27232
rect 32692 27172 32696 27228
rect 32696 27172 32752 27228
rect 32752 27172 32756 27228
rect 32692 27168 32756 27172
rect 32772 27228 32836 27232
rect 32772 27172 32776 27228
rect 32776 27172 32832 27228
rect 32832 27172 32836 27228
rect 32772 27168 32836 27172
rect 32852 27228 32916 27232
rect 32852 27172 32856 27228
rect 32856 27172 32912 27228
rect 32912 27172 32916 27228
rect 32852 27168 32916 27172
rect 37612 27228 37676 27232
rect 37612 27172 37616 27228
rect 37616 27172 37672 27228
rect 37672 27172 37676 27228
rect 37612 27168 37676 27172
rect 37692 27228 37756 27232
rect 37692 27172 37696 27228
rect 37696 27172 37752 27228
rect 37752 27172 37756 27228
rect 37692 27168 37756 27172
rect 37772 27228 37836 27232
rect 37772 27172 37776 27228
rect 37776 27172 37832 27228
rect 37832 27172 37836 27228
rect 37772 27168 37836 27172
rect 37852 27228 37916 27232
rect 37852 27172 37856 27228
rect 37856 27172 37912 27228
rect 37912 27172 37916 27228
rect 37852 27168 37916 27172
rect 1952 26684 2016 26688
rect 1952 26628 1956 26684
rect 1956 26628 2012 26684
rect 2012 26628 2016 26684
rect 1952 26624 2016 26628
rect 2032 26684 2096 26688
rect 2032 26628 2036 26684
rect 2036 26628 2092 26684
rect 2092 26628 2096 26684
rect 2032 26624 2096 26628
rect 2112 26684 2176 26688
rect 2112 26628 2116 26684
rect 2116 26628 2172 26684
rect 2172 26628 2176 26684
rect 2112 26624 2176 26628
rect 2192 26684 2256 26688
rect 2192 26628 2196 26684
rect 2196 26628 2252 26684
rect 2252 26628 2256 26684
rect 2192 26624 2256 26628
rect 6952 26684 7016 26688
rect 6952 26628 6956 26684
rect 6956 26628 7012 26684
rect 7012 26628 7016 26684
rect 6952 26624 7016 26628
rect 7032 26684 7096 26688
rect 7032 26628 7036 26684
rect 7036 26628 7092 26684
rect 7092 26628 7096 26684
rect 7032 26624 7096 26628
rect 7112 26684 7176 26688
rect 7112 26628 7116 26684
rect 7116 26628 7172 26684
rect 7172 26628 7176 26684
rect 7112 26624 7176 26628
rect 7192 26684 7256 26688
rect 7192 26628 7196 26684
rect 7196 26628 7252 26684
rect 7252 26628 7256 26684
rect 7192 26624 7256 26628
rect 11952 26684 12016 26688
rect 11952 26628 11956 26684
rect 11956 26628 12012 26684
rect 12012 26628 12016 26684
rect 11952 26624 12016 26628
rect 12032 26684 12096 26688
rect 12032 26628 12036 26684
rect 12036 26628 12092 26684
rect 12092 26628 12096 26684
rect 12032 26624 12096 26628
rect 12112 26684 12176 26688
rect 12112 26628 12116 26684
rect 12116 26628 12172 26684
rect 12172 26628 12176 26684
rect 12112 26624 12176 26628
rect 12192 26684 12256 26688
rect 12192 26628 12196 26684
rect 12196 26628 12252 26684
rect 12252 26628 12256 26684
rect 12192 26624 12256 26628
rect 16952 26684 17016 26688
rect 16952 26628 16956 26684
rect 16956 26628 17012 26684
rect 17012 26628 17016 26684
rect 16952 26624 17016 26628
rect 17032 26684 17096 26688
rect 17032 26628 17036 26684
rect 17036 26628 17092 26684
rect 17092 26628 17096 26684
rect 17032 26624 17096 26628
rect 17112 26684 17176 26688
rect 17112 26628 17116 26684
rect 17116 26628 17172 26684
rect 17172 26628 17176 26684
rect 17112 26624 17176 26628
rect 17192 26684 17256 26688
rect 17192 26628 17196 26684
rect 17196 26628 17252 26684
rect 17252 26628 17256 26684
rect 17192 26624 17256 26628
rect 21952 26684 22016 26688
rect 21952 26628 21956 26684
rect 21956 26628 22012 26684
rect 22012 26628 22016 26684
rect 21952 26624 22016 26628
rect 22032 26684 22096 26688
rect 22032 26628 22036 26684
rect 22036 26628 22092 26684
rect 22092 26628 22096 26684
rect 22032 26624 22096 26628
rect 22112 26684 22176 26688
rect 22112 26628 22116 26684
rect 22116 26628 22172 26684
rect 22172 26628 22176 26684
rect 22112 26624 22176 26628
rect 22192 26684 22256 26688
rect 22192 26628 22196 26684
rect 22196 26628 22252 26684
rect 22252 26628 22256 26684
rect 22192 26624 22256 26628
rect 26952 26684 27016 26688
rect 26952 26628 26956 26684
rect 26956 26628 27012 26684
rect 27012 26628 27016 26684
rect 26952 26624 27016 26628
rect 27032 26684 27096 26688
rect 27032 26628 27036 26684
rect 27036 26628 27092 26684
rect 27092 26628 27096 26684
rect 27032 26624 27096 26628
rect 27112 26684 27176 26688
rect 27112 26628 27116 26684
rect 27116 26628 27172 26684
rect 27172 26628 27176 26684
rect 27112 26624 27176 26628
rect 27192 26684 27256 26688
rect 27192 26628 27196 26684
rect 27196 26628 27252 26684
rect 27252 26628 27256 26684
rect 27192 26624 27256 26628
rect 31952 26684 32016 26688
rect 31952 26628 31956 26684
rect 31956 26628 32012 26684
rect 32012 26628 32016 26684
rect 31952 26624 32016 26628
rect 32032 26684 32096 26688
rect 32032 26628 32036 26684
rect 32036 26628 32092 26684
rect 32092 26628 32096 26684
rect 32032 26624 32096 26628
rect 32112 26684 32176 26688
rect 32112 26628 32116 26684
rect 32116 26628 32172 26684
rect 32172 26628 32176 26684
rect 32112 26624 32176 26628
rect 32192 26684 32256 26688
rect 32192 26628 32196 26684
rect 32196 26628 32252 26684
rect 32252 26628 32256 26684
rect 32192 26624 32256 26628
rect 36952 26684 37016 26688
rect 36952 26628 36956 26684
rect 36956 26628 37012 26684
rect 37012 26628 37016 26684
rect 36952 26624 37016 26628
rect 37032 26684 37096 26688
rect 37032 26628 37036 26684
rect 37036 26628 37092 26684
rect 37092 26628 37096 26684
rect 37032 26624 37096 26628
rect 37112 26684 37176 26688
rect 37112 26628 37116 26684
rect 37116 26628 37172 26684
rect 37172 26628 37176 26684
rect 37112 26624 37176 26628
rect 37192 26684 37256 26688
rect 37192 26628 37196 26684
rect 37196 26628 37252 26684
rect 37252 26628 37256 26684
rect 37192 26624 37256 26628
rect 2612 26140 2676 26144
rect 2612 26084 2616 26140
rect 2616 26084 2672 26140
rect 2672 26084 2676 26140
rect 2612 26080 2676 26084
rect 2692 26140 2756 26144
rect 2692 26084 2696 26140
rect 2696 26084 2752 26140
rect 2752 26084 2756 26140
rect 2692 26080 2756 26084
rect 2772 26140 2836 26144
rect 2772 26084 2776 26140
rect 2776 26084 2832 26140
rect 2832 26084 2836 26140
rect 2772 26080 2836 26084
rect 2852 26140 2916 26144
rect 2852 26084 2856 26140
rect 2856 26084 2912 26140
rect 2912 26084 2916 26140
rect 2852 26080 2916 26084
rect 7612 26140 7676 26144
rect 7612 26084 7616 26140
rect 7616 26084 7672 26140
rect 7672 26084 7676 26140
rect 7612 26080 7676 26084
rect 7692 26140 7756 26144
rect 7692 26084 7696 26140
rect 7696 26084 7752 26140
rect 7752 26084 7756 26140
rect 7692 26080 7756 26084
rect 7772 26140 7836 26144
rect 7772 26084 7776 26140
rect 7776 26084 7832 26140
rect 7832 26084 7836 26140
rect 7772 26080 7836 26084
rect 7852 26140 7916 26144
rect 7852 26084 7856 26140
rect 7856 26084 7912 26140
rect 7912 26084 7916 26140
rect 7852 26080 7916 26084
rect 12612 26140 12676 26144
rect 12612 26084 12616 26140
rect 12616 26084 12672 26140
rect 12672 26084 12676 26140
rect 12612 26080 12676 26084
rect 12692 26140 12756 26144
rect 12692 26084 12696 26140
rect 12696 26084 12752 26140
rect 12752 26084 12756 26140
rect 12692 26080 12756 26084
rect 12772 26140 12836 26144
rect 12772 26084 12776 26140
rect 12776 26084 12832 26140
rect 12832 26084 12836 26140
rect 12772 26080 12836 26084
rect 12852 26140 12916 26144
rect 12852 26084 12856 26140
rect 12856 26084 12912 26140
rect 12912 26084 12916 26140
rect 12852 26080 12916 26084
rect 17612 26140 17676 26144
rect 17612 26084 17616 26140
rect 17616 26084 17672 26140
rect 17672 26084 17676 26140
rect 17612 26080 17676 26084
rect 17692 26140 17756 26144
rect 17692 26084 17696 26140
rect 17696 26084 17752 26140
rect 17752 26084 17756 26140
rect 17692 26080 17756 26084
rect 17772 26140 17836 26144
rect 17772 26084 17776 26140
rect 17776 26084 17832 26140
rect 17832 26084 17836 26140
rect 17772 26080 17836 26084
rect 17852 26140 17916 26144
rect 17852 26084 17856 26140
rect 17856 26084 17912 26140
rect 17912 26084 17916 26140
rect 17852 26080 17916 26084
rect 22612 26140 22676 26144
rect 22612 26084 22616 26140
rect 22616 26084 22672 26140
rect 22672 26084 22676 26140
rect 22612 26080 22676 26084
rect 22692 26140 22756 26144
rect 22692 26084 22696 26140
rect 22696 26084 22752 26140
rect 22752 26084 22756 26140
rect 22692 26080 22756 26084
rect 22772 26140 22836 26144
rect 22772 26084 22776 26140
rect 22776 26084 22832 26140
rect 22832 26084 22836 26140
rect 22772 26080 22836 26084
rect 22852 26140 22916 26144
rect 22852 26084 22856 26140
rect 22856 26084 22912 26140
rect 22912 26084 22916 26140
rect 22852 26080 22916 26084
rect 27612 26140 27676 26144
rect 27612 26084 27616 26140
rect 27616 26084 27672 26140
rect 27672 26084 27676 26140
rect 27612 26080 27676 26084
rect 27692 26140 27756 26144
rect 27692 26084 27696 26140
rect 27696 26084 27752 26140
rect 27752 26084 27756 26140
rect 27692 26080 27756 26084
rect 27772 26140 27836 26144
rect 27772 26084 27776 26140
rect 27776 26084 27832 26140
rect 27832 26084 27836 26140
rect 27772 26080 27836 26084
rect 27852 26140 27916 26144
rect 27852 26084 27856 26140
rect 27856 26084 27912 26140
rect 27912 26084 27916 26140
rect 27852 26080 27916 26084
rect 32612 26140 32676 26144
rect 32612 26084 32616 26140
rect 32616 26084 32672 26140
rect 32672 26084 32676 26140
rect 32612 26080 32676 26084
rect 32692 26140 32756 26144
rect 32692 26084 32696 26140
rect 32696 26084 32752 26140
rect 32752 26084 32756 26140
rect 32692 26080 32756 26084
rect 32772 26140 32836 26144
rect 32772 26084 32776 26140
rect 32776 26084 32832 26140
rect 32832 26084 32836 26140
rect 32772 26080 32836 26084
rect 32852 26140 32916 26144
rect 32852 26084 32856 26140
rect 32856 26084 32912 26140
rect 32912 26084 32916 26140
rect 32852 26080 32916 26084
rect 37612 26140 37676 26144
rect 37612 26084 37616 26140
rect 37616 26084 37672 26140
rect 37672 26084 37676 26140
rect 37612 26080 37676 26084
rect 37692 26140 37756 26144
rect 37692 26084 37696 26140
rect 37696 26084 37752 26140
rect 37752 26084 37756 26140
rect 37692 26080 37756 26084
rect 37772 26140 37836 26144
rect 37772 26084 37776 26140
rect 37776 26084 37832 26140
rect 37832 26084 37836 26140
rect 37772 26080 37836 26084
rect 37852 26140 37916 26144
rect 37852 26084 37856 26140
rect 37856 26084 37912 26140
rect 37912 26084 37916 26140
rect 37852 26080 37916 26084
rect 1952 25596 2016 25600
rect 1952 25540 1956 25596
rect 1956 25540 2012 25596
rect 2012 25540 2016 25596
rect 1952 25536 2016 25540
rect 2032 25596 2096 25600
rect 2032 25540 2036 25596
rect 2036 25540 2092 25596
rect 2092 25540 2096 25596
rect 2032 25536 2096 25540
rect 2112 25596 2176 25600
rect 2112 25540 2116 25596
rect 2116 25540 2172 25596
rect 2172 25540 2176 25596
rect 2112 25536 2176 25540
rect 2192 25596 2256 25600
rect 2192 25540 2196 25596
rect 2196 25540 2252 25596
rect 2252 25540 2256 25596
rect 2192 25536 2256 25540
rect 6952 25596 7016 25600
rect 6952 25540 6956 25596
rect 6956 25540 7012 25596
rect 7012 25540 7016 25596
rect 6952 25536 7016 25540
rect 7032 25596 7096 25600
rect 7032 25540 7036 25596
rect 7036 25540 7092 25596
rect 7092 25540 7096 25596
rect 7032 25536 7096 25540
rect 7112 25596 7176 25600
rect 7112 25540 7116 25596
rect 7116 25540 7172 25596
rect 7172 25540 7176 25596
rect 7112 25536 7176 25540
rect 7192 25596 7256 25600
rect 7192 25540 7196 25596
rect 7196 25540 7252 25596
rect 7252 25540 7256 25596
rect 7192 25536 7256 25540
rect 11952 25596 12016 25600
rect 11952 25540 11956 25596
rect 11956 25540 12012 25596
rect 12012 25540 12016 25596
rect 11952 25536 12016 25540
rect 12032 25596 12096 25600
rect 12032 25540 12036 25596
rect 12036 25540 12092 25596
rect 12092 25540 12096 25596
rect 12032 25536 12096 25540
rect 12112 25596 12176 25600
rect 12112 25540 12116 25596
rect 12116 25540 12172 25596
rect 12172 25540 12176 25596
rect 12112 25536 12176 25540
rect 12192 25596 12256 25600
rect 12192 25540 12196 25596
rect 12196 25540 12252 25596
rect 12252 25540 12256 25596
rect 12192 25536 12256 25540
rect 16952 25596 17016 25600
rect 16952 25540 16956 25596
rect 16956 25540 17012 25596
rect 17012 25540 17016 25596
rect 16952 25536 17016 25540
rect 17032 25596 17096 25600
rect 17032 25540 17036 25596
rect 17036 25540 17092 25596
rect 17092 25540 17096 25596
rect 17032 25536 17096 25540
rect 17112 25596 17176 25600
rect 17112 25540 17116 25596
rect 17116 25540 17172 25596
rect 17172 25540 17176 25596
rect 17112 25536 17176 25540
rect 17192 25596 17256 25600
rect 17192 25540 17196 25596
rect 17196 25540 17252 25596
rect 17252 25540 17256 25596
rect 17192 25536 17256 25540
rect 21952 25596 22016 25600
rect 21952 25540 21956 25596
rect 21956 25540 22012 25596
rect 22012 25540 22016 25596
rect 21952 25536 22016 25540
rect 22032 25596 22096 25600
rect 22032 25540 22036 25596
rect 22036 25540 22092 25596
rect 22092 25540 22096 25596
rect 22032 25536 22096 25540
rect 22112 25596 22176 25600
rect 22112 25540 22116 25596
rect 22116 25540 22172 25596
rect 22172 25540 22176 25596
rect 22112 25536 22176 25540
rect 22192 25596 22256 25600
rect 22192 25540 22196 25596
rect 22196 25540 22252 25596
rect 22252 25540 22256 25596
rect 22192 25536 22256 25540
rect 26952 25596 27016 25600
rect 26952 25540 26956 25596
rect 26956 25540 27012 25596
rect 27012 25540 27016 25596
rect 26952 25536 27016 25540
rect 27032 25596 27096 25600
rect 27032 25540 27036 25596
rect 27036 25540 27092 25596
rect 27092 25540 27096 25596
rect 27032 25536 27096 25540
rect 27112 25596 27176 25600
rect 27112 25540 27116 25596
rect 27116 25540 27172 25596
rect 27172 25540 27176 25596
rect 27112 25536 27176 25540
rect 27192 25596 27256 25600
rect 27192 25540 27196 25596
rect 27196 25540 27252 25596
rect 27252 25540 27256 25596
rect 27192 25536 27256 25540
rect 31952 25596 32016 25600
rect 31952 25540 31956 25596
rect 31956 25540 32012 25596
rect 32012 25540 32016 25596
rect 31952 25536 32016 25540
rect 32032 25596 32096 25600
rect 32032 25540 32036 25596
rect 32036 25540 32092 25596
rect 32092 25540 32096 25596
rect 32032 25536 32096 25540
rect 32112 25596 32176 25600
rect 32112 25540 32116 25596
rect 32116 25540 32172 25596
rect 32172 25540 32176 25596
rect 32112 25536 32176 25540
rect 32192 25596 32256 25600
rect 32192 25540 32196 25596
rect 32196 25540 32252 25596
rect 32252 25540 32256 25596
rect 32192 25536 32256 25540
rect 36952 25596 37016 25600
rect 36952 25540 36956 25596
rect 36956 25540 37012 25596
rect 37012 25540 37016 25596
rect 36952 25536 37016 25540
rect 37032 25596 37096 25600
rect 37032 25540 37036 25596
rect 37036 25540 37092 25596
rect 37092 25540 37096 25596
rect 37032 25536 37096 25540
rect 37112 25596 37176 25600
rect 37112 25540 37116 25596
rect 37116 25540 37172 25596
rect 37172 25540 37176 25596
rect 37112 25536 37176 25540
rect 37192 25596 37256 25600
rect 37192 25540 37196 25596
rect 37196 25540 37252 25596
rect 37252 25540 37256 25596
rect 37192 25536 37256 25540
rect 2612 25052 2676 25056
rect 2612 24996 2616 25052
rect 2616 24996 2672 25052
rect 2672 24996 2676 25052
rect 2612 24992 2676 24996
rect 2692 25052 2756 25056
rect 2692 24996 2696 25052
rect 2696 24996 2752 25052
rect 2752 24996 2756 25052
rect 2692 24992 2756 24996
rect 2772 25052 2836 25056
rect 2772 24996 2776 25052
rect 2776 24996 2832 25052
rect 2832 24996 2836 25052
rect 2772 24992 2836 24996
rect 2852 25052 2916 25056
rect 2852 24996 2856 25052
rect 2856 24996 2912 25052
rect 2912 24996 2916 25052
rect 2852 24992 2916 24996
rect 7612 25052 7676 25056
rect 7612 24996 7616 25052
rect 7616 24996 7672 25052
rect 7672 24996 7676 25052
rect 7612 24992 7676 24996
rect 7692 25052 7756 25056
rect 7692 24996 7696 25052
rect 7696 24996 7752 25052
rect 7752 24996 7756 25052
rect 7692 24992 7756 24996
rect 7772 25052 7836 25056
rect 7772 24996 7776 25052
rect 7776 24996 7832 25052
rect 7832 24996 7836 25052
rect 7772 24992 7836 24996
rect 7852 25052 7916 25056
rect 7852 24996 7856 25052
rect 7856 24996 7912 25052
rect 7912 24996 7916 25052
rect 7852 24992 7916 24996
rect 12612 25052 12676 25056
rect 12612 24996 12616 25052
rect 12616 24996 12672 25052
rect 12672 24996 12676 25052
rect 12612 24992 12676 24996
rect 12692 25052 12756 25056
rect 12692 24996 12696 25052
rect 12696 24996 12752 25052
rect 12752 24996 12756 25052
rect 12692 24992 12756 24996
rect 12772 25052 12836 25056
rect 12772 24996 12776 25052
rect 12776 24996 12832 25052
rect 12832 24996 12836 25052
rect 12772 24992 12836 24996
rect 12852 25052 12916 25056
rect 12852 24996 12856 25052
rect 12856 24996 12912 25052
rect 12912 24996 12916 25052
rect 12852 24992 12916 24996
rect 17612 25052 17676 25056
rect 17612 24996 17616 25052
rect 17616 24996 17672 25052
rect 17672 24996 17676 25052
rect 17612 24992 17676 24996
rect 17692 25052 17756 25056
rect 17692 24996 17696 25052
rect 17696 24996 17752 25052
rect 17752 24996 17756 25052
rect 17692 24992 17756 24996
rect 17772 25052 17836 25056
rect 17772 24996 17776 25052
rect 17776 24996 17832 25052
rect 17832 24996 17836 25052
rect 17772 24992 17836 24996
rect 17852 25052 17916 25056
rect 17852 24996 17856 25052
rect 17856 24996 17912 25052
rect 17912 24996 17916 25052
rect 17852 24992 17916 24996
rect 22612 25052 22676 25056
rect 22612 24996 22616 25052
rect 22616 24996 22672 25052
rect 22672 24996 22676 25052
rect 22612 24992 22676 24996
rect 22692 25052 22756 25056
rect 22692 24996 22696 25052
rect 22696 24996 22752 25052
rect 22752 24996 22756 25052
rect 22692 24992 22756 24996
rect 22772 25052 22836 25056
rect 22772 24996 22776 25052
rect 22776 24996 22832 25052
rect 22832 24996 22836 25052
rect 22772 24992 22836 24996
rect 22852 25052 22916 25056
rect 22852 24996 22856 25052
rect 22856 24996 22912 25052
rect 22912 24996 22916 25052
rect 22852 24992 22916 24996
rect 27612 25052 27676 25056
rect 27612 24996 27616 25052
rect 27616 24996 27672 25052
rect 27672 24996 27676 25052
rect 27612 24992 27676 24996
rect 27692 25052 27756 25056
rect 27692 24996 27696 25052
rect 27696 24996 27752 25052
rect 27752 24996 27756 25052
rect 27692 24992 27756 24996
rect 27772 25052 27836 25056
rect 27772 24996 27776 25052
rect 27776 24996 27832 25052
rect 27832 24996 27836 25052
rect 27772 24992 27836 24996
rect 27852 25052 27916 25056
rect 27852 24996 27856 25052
rect 27856 24996 27912 25052
rect 27912 24996 27916 25052
rect 27852 24992 27916 24996
rect 32612 25052 32676 25056
rect 32612 24996 32616 25052
rect 32616 24996 32672 25052
rect 32672 24996 32676 25052
rect 32612 24992 32676 24996
rect 32692 25052 32756 25056
rect 32692 24996 32696 25052
rect 32696 24996 32752 25052
rect 32752 24996 32756 25052
rect 32692 24992 32756 24996
rect 32772 25052 32836 25056
rect 32772 24996 32776 25052
rect 32776 24996 32832 25052
rect 32832 24996 32836 25052
rect 32772 24992 32836 24996
rect 32852 25052 32916 25056
rect 32852 24996 32856 25052
rect 32856 24996 32912 25052
rect 32912 24996 32916 25052
rect 32852 24992 32916 24996
rect 37612 25052 37676 25056
rect 37612 24996 37616 25052
rect 37616 24996 37672 25052
rect 37672 24996 37676 25052
rect 37612 24992 37676 24996
rect 37692 25052 37756 25056
rect 37692 24996 37696 25052
rect 37696 24996 37752 25052
rect 37752 24996 37756 25052
rect 37692 24992 37756 24996
rect 37772 25052 37836 25056
rect 37772 24996 37776 25052
rect 37776 24996 37832 25052
rect 37832 24996 37836 25052
rect 37772 24992 37836 24996
rect 37852 25052 37916 25056
rect 37852 24996 37856 25052
rect 37856 24996 37912 25052
rect 37912 24996 37916 25052
rect 37852 24992 37916 24996
rect 1952 24508 2016 24512
rect 1952 24452 1956 24508
rect 1956 24452 2012 24508
rect 2012 24452 2016 24508
rect 1952 24448 2016 24452
rect 2032 24508 2096 24512
rect 2032 24452 2036 24508
rect 2036 24452 2092 24508
rect 2092 24452 2096 24508
rect 2032 24448 2096 24452
rect 2112 24508 2176 24512
rect 2112 24452 2116 24508
rect 2116 24452 2172 24508
rect 2172 24452 2176 24508
rect 2112 24448 2176 24452
rect 2192 24508 2256 24512
rect 2192 24452 2196 24508
rect 2196 24452 2252 24508
rect 2252 24452 2256 24508
rect 2192 24448 2256 24452
rect 6952 24508 7016 24512
rect 6952 24452 6956 24508
rect 6956 24452 7012 24508
rect 7012 24452 7016 24508
rect 6952 24448 7016 24452
rect 7032 24508 7096 24512
rect 7032 24452 7036 24508
rect 7036 24452 7092 24508
rect 7092 24452 7096 24508
rect 7032 24448 7096 24452
rect 7112 24508 7176 24512
rect 7112 24452 7116 24508
rect 7116 24452 7172 24508
rect 7172 24452 7176 24508
rect 7112 24448 7176 24452
rect 7192 24508 7256 24512
rect 7192 24452 7196 24508
rect 7196 24452 7252 24508
rect 7252 24452 7256 24508
rect 7192 24448 7256 24452
rect 11952 24508 12016 24512
rect 11952 24452 11956 24508
rect 11956 24452 12012 24508
rect 12012 24452 12016 24508
rect 11952 24448 12016 24452
rect 12032 24508 12096 24512
rect 12032 24452 12036 24508
rect 12036 24452 12092 24508
rect 12092 24452 12096 24508
rect 12032 24448 12096 24452
rect 12112 24508 12176 24512
rect 12112 24452 12116 24508
rect 12116 24452 12172 24508
rect 12172 24452 12176 24508
rect 12112 24448 12176 24452
rect 12192 24508 12256 24512
rect 12192 24452 12196 24508
rect 12196 24452 12252 24508
rect 12252 24452 12256 24508
rect 12192 24448 12256 24452
rect 16952 24508 17016 24512
rect 16952 24452 16956 24508
rect 16956 24452 17012 24508
rect 17012 24452 17016 24508
rect 16952 24448 17016 24452
rect 17032 24508 17096 24512
rect 17032 24452 17036 24508
rect 17036 24452 17092 24508
rect 17092 24452 17096 24508
rect 17032 24448 17096 24452
rect 17112 24508 17176 24512
rect 17112 24452 17116 24508
rect 17116 24452 17172 24508
rect 17172 24452 17176 24508
rect 17112 24448 17176 24452
rect 17192 24508 17256 24512
rect 17192 24452 17196 24508
rect 17196 24452 17252 24508
rect 17252 24452 17256 24508
rect 17192 24448 17256 24452
rect 21952 24508 22016 24512
rect 21952 24452 21956 24508
rect 21956 24452 22012 24508
rect 22012 24452 22016 24508
rect 21952 24448 22016 24452
rect 22032 24508 22096 24512
rect 22032 24452 22036 24508
rect 22036 24452 22092 24508
rect 22092 24452 22096 24508
rect 22032 24448 22096 24452
rect 22112 24508 22176 24512
rect 22112 24452 22116 24508
rect 22116 24452 22172 24508
rect 22172 24452 22176 24508
rect 22112 24448 22176 24452
rect 22192 24508 22256 24512
rect 22192 24452 22196 24508
rect 22196 24452 22252 24508
rect 22252 24452 22256 24508
rect 22192 24448 22256 24452
rect 26952 24508 27016 24512
rect 26952 24452 26956 24508
rect 26956 24452 27012 24508
rect 27012 24452 27016 24508
rect 26952 24448 27016 24452
rect 27032 24508 27096 24512
rect 27032 24452 27036 24508
rect 27036 24452 27092 24508
rect 27092 24452 27096 24508
rect 27032 24448 27096 24452
rect 27112 24508 27176 24512
rect 27112 24452 27116 24508
rect 27116 24452 27172 24508
rect 27172 24452 27176 24508
rect 27112 24448 27176 24452
rect 27192 24508 27256 24512
rect 27192 24452 27196 24508
rect 27196 24452 27252 24508
rect 27252 24452 27256 24508
rect 27192 24448 27256 24452
rect 31952 24508 32016 24512
rect 31952 24452 31956 24508
rect 31956 24452 32012 24508
rect 32012 24452 32016 24508
rect 31952 24448 32016 24452
rect 32032 24508 32096 24512
rect 32032 24452 32036 24508
rect 32036 24452 32092 24508
rect 32092 24452 32096 24508
rect 32032 24448 32096 24452
rect 32112 24508 32176 24512
rect 32112 24452 32116 24508
rect 32116 24452 32172 24508
rect 32172 24452 32176 24508
rect 32112 24448 32176 24452
rect 32192 24508 32256 24512
rect 32192 24452 32196 24508
rect 32196 24452 32252 24508
rect 32252 24452 32256 24508
rect 32192 24448 32256 24452
rect 36952 24508 37016 24512
rect 36952 24452 36956 24508
rect 36956 24452 37012 24508
rect 37012 24452 37016 24508
rect 36952 24448 37016 24452
rect 37032 24508 37096 24512
rect 37032 24452 37036 24508
rect 37036 24452 37092 24508
rect 37092 24452 37096 24508
rect 37032 24448 37096 24452
rect 37112 24508 37176 24512
rect 37112 24452 37116 24508
rect 37116 24452 37172 24508
rect 37172 24452 37176 24508
rect 37112 24448 37176 24452
rect 37192 24508 37256 24512
rect 37192 24452 37196 24508
rect 37196 24452 37252 24508
rect 37252 24452 37256 24508
rect 37192 24448 37256 24452
rect 2612 23964 2676 23968
rect 2612 23908 2616 23964
rect 2616 23908 2672 23964
rect 2672 23908 2676 23964
rect 2612 23904 2676 23908
rect 2692 23964 2756 23968
rect 2692 23908 2696 23964
rect 2696 23908 2752 23964
rect 2752 23908 2756 23964
rect 2692 23904 2756 23908
rect 2772 23964 2836 23968
rect 2772 23908 2776 23964
rect 2776 23908 2832 23964
rect 2832 23908 2836 23964
rect 2772 23904 2836 23908
rect 2852 23964 2916 23968
rect 2852 23908 2856 23964
rect 2856 23908 2912 23964
rect 2912 23908 2916 23964
rect 2852 23904 2916 23908
rect 7612 23964 7676 23968
rect 7612 23908 7616 23964
rect 7616 23908 7672 23964
rect 7672 23908 7676 23964
rect 7612 23904 7676 23908
rect 7692 23964 7756 23968
rect 7692 23908 7696 23964
rect 7696 23908 7752 23964
rect 7752 23908 7756 23964
rect 7692 23904 7756 23908
rect 7772 23964 7836 23968
rect 7772 23908 7776 23964
rect 7776 23908 7832 23964
rect 7832 23908 7836 23964
rect 7772 23904 7836 23908
rect 7852 23964 7916 23968
rect 7852 23908 7856 23964
rect 7856 23908 7912 23964
rect 7912 23908 7916 23964
rect 7852 23904 7916 23908
rect 12612 23964 12676 23968
rect 12612 23908 12616 23964
rect 12616 23908 12672 23964
rect 12672 23908 12676 23964
rect 12612 23904 12676 23908
rect 12692 23964 12756 23968
rect 12692 23908 12696 23964
rect 12696 23908 12752 23964
rect 12752 23908 12756 23964
rect 12692 23904 12756 23908
rect 12772 23964 12836 23968
rect 12772 23908 12776 23964
rect 12776 23908 12832 23964
rect 12832 23908 12836 23964
rect 12772 23904 12836 23908
rect 12852 23964 12916 23968
rect 12852 23908 12856 23964
rect 12856 23908 12912 23964
rect 12912 23908 12916 23964
rect 12852 23904 12916 23908
rect 17612 23964 17676 23968
rect 17612 23908 17616 23964
rect 17616 23908 17672 23964
rect 17672 23908 17676 23964
rect 17612 23904 17676 23908
rect 17692 23964 17756 23968
rect 17692 23908 17696 23964
rect 17696 23908 17752 23964
rect 17752 23908 17756 23964
rect 17692 23904 17756 23908
rect 17772 23964 17836 23968
rect 17772 23908 17776 23964
rect 17776 23908 17832 23964
rect 17832 23908 17836 23964
rect 17772 23904 17836 23908
rect 17852 23964 17916 23968
rect 17852 23908 17856 23964
rect 17856 23908 17912 23964
rect 17912 23908 17916 23964
rect 17852 23904 17916 23908
rect 22612 23964 22676 23968
rect 22612 23908 22616 23964
rect 22616 23908 22672 23964
rect 22672 23908 22676 23964
rect 22612 23904 22676 23908
rect 22692 23964 22756 23968
rect 22692 23908 22696 23964
rect 22696 23908 22752 23964
rect 22752 23908 22756 23964
rect 22692 23904 22756 23908
rect 22772 23964 22836 23968
rect 22772 23908 22776 23964
rect 22776 23908 22832 23964
rect 22832 23908 22836 23964
rect 22772 23904 22836 23908
rect 22852 23964 22916 23968
rect 22852 23908 22856 23964
rect 22856 23908 22912 23964
rect 22912 23908 22916 23964
rect 22852 23904 22916 23908
rect 27612 23964 27676 23968
rect 27612 23908 27616 23964
rect 27616 23908 27672 23964
rect 27672 23908 27676 23964
rect 27612 23904 27676 23908
rect 27692 23964 27756 23968
rect 27692 23908 27696 23964
rect 27696 23908 27752 23964
rect 27752 23908 27756 23964
rect 27692 23904 27756 23908
rect 27772 23964 27836 23968
rect 27772 23908 27776 23964
rect 27776 23908 27832 23964
rect 27832 23908 27836 23964
rect 27772 23904 27836 23908
rect 27852 23964 27916 23968
rect 27852 23908 27856 23964
rect 27856 23908 27912 23964
rect 27912 23908 27916 23964
rect 27852 23904 27916 23908
rect 32612 23964 32676 23968
rect 32612 23908 32616 23964
rect 32616 23908 32672 23964
rect 32672 23908 32676 23964
rect 32612 23904 32676 23908
rect 32692 23964 32756 23968
rect 32692 23908 32696 23964
rect 32696 23908 32752 23964
rect 32752 23908 32756 23964
rect 32692 23904 32756 23908
rect 32772 23964 32836 23968
rect 32772 23908 32776 23964
rect 32776 23908 32832 23964
rect 32832 23908 32836 23964
rect 32772 23904 32836 23908
rect 32852 23964 32916 23968
rect 32852 23908 32856 23964
rect 32856 23908 32912 23964
rect 32912 23908 32916 23964
rect 32852 23904 32916 23908
rect 37612 23964 37676 23968
rect 37612 23908 37616 23964
rect 37616 23908 37672 23964
rect 37672 23908 37676 23964
rect 37612 23904 37676 23908
rect 37692 23964 37756 23968
rect 37692 23908 37696 23964
rect 37696 23908 37752 23964
rect 37752 23908 37756 23964
rect 37692 23904 37756 23908
rect 37772 23964 37836 23968
rect 37772 23908 37776 23964
rect 37776 23908 37832 23964
rect 37832 23908 37836 23964
rect 37772 23904 37836 23908
rect 37852 23964 37916 23968
rect 37852 23908 37856 23964
rect 37856 23908 37912 23964
rect 37912 23908 37916 23964
rect 37852 23904 37916 23908
rect 1952 23420 2016 23424
rect 1952 23364 1956 23420
rect 1956 23364 2012 23420
rect 2012 23364 2016 23420
rect 1952 23360 2016 23364
rect 2032 23420 2096 23424
rect 2032 23364 2036 23420
rect 2036 23364 2092 23420
rect 2092 23364 2096 23420
rect 2032 23360 2096 23364
rect 2112 23420 2176 23424
rect 2112 23364 2116 23420
rect 2116 23364 2172 23420
rect 2172 23364 2176 23420
rect 2112 23360 2176 23364
rect 2192 23420 2256 23424
rect 2192 23364 2196 23420
rect 2196 23364 2252 23420
rect 2252 23364 2256 23420
rect 2192 23360 2256 23364
rect 6952 23420 7016 23424
rect 6952 23364 6956 23420
rect 6956 23364 7012 23420
rect 7012 23364 7016 23420
rect 6952 23360 7016 23364
rect 7032 23420 7096 23424
rect 7032 23364 7036 23420
rect 7036 23364 7092 23420
rect 7092 23364 7096 23420
rect 7032 23360 7096 23364
rect 7112 23420 7176 23424
rect 7112 23364 7116 23420
rect 7116 23364 7172 23420
rect 7172 23364 7176 23420
rect 7112 23360 7176 23364
rect 7192 23420 7256 23424
rect 7192 23364 7196 23420
rect 7196 23364 7252 23420
rect 7252 23364 7256 23420
rect 7192 23360 7256 23364
rect 11952 23420 12016 23424
rect 11952 23364 11956 23420
rect 11956 23364 12012 23420
rect 12012 23364 12016 23420
rect 11952 23360 12016 23364
rect 12032 23420 12096 23424
rect 12032 23364 12036 23420
rect 12036 23364 12092 23420
rect 12092 23364 12096 23420
rect 12032 23360 12096 23364
rect 12112 23420 12176 23424
rect 12112 23364 12116 23420
rect 12116 23364 12172 23420
rect 12172 23364 12176 23420
rect 12112 23360 12176 23364
rect 12192 23420 12256 23424
rect 12192 23364 12196 23420
rect 12196 23364 12252 23420
rect 12252 23364 12256 23420
rect 12192 23360 12256 23364
rect 16952 23420 17016 23424
rect 16952 23364 16956 23420
rect 16956 23364 17012 23420
rect 17012 23364 17016 23420
rect 16952 23360 17016 23364
rect 17032 23420 17096 23424
rect 17032 23364 17036 23420
rect 17036 23364 17092 23420
rect 17092 23364 17096 23420
rect 17032 23360 17096 23364
rect 17112 23420 17176 23424
rect 17112 23364 17116 23420
rect 17116 23364 17172 23420
rect 17172 23364 17176 23420
rect 17112 23360 17176 23364
rect 17192 23420 17256 23424
rect 17192 23364 17196 23420
rect 17196 23364 17252 23420
rect 17252 23364 17256 23420
rect 17192 23360 17256 23364
rect 21952 23420 22016 23424
rect 21952 23364 21956 23420
rect 21956 23364 22012 23420
rect 22012 23364 22016 23420
rect 21952 23360 22016 23364
rect 22032 23420 22096 23424
rect 22032 23364 22036 23420
rect 22036 23364 22092 23420
rect 22092 23364 22096 23420
rect 22032 23360 22096 23364
rect 22112 23420 22176 23424
rect 22112 23364 22116 23420
rect 22116 23364 22172 23420
rect 22172 23364 22176 23420
rect 22112 23360 22176 23364
rect 22192 23420 22256 23424
rect 22192 23364 22196 23420
rect 22196 23364 22252 23420
rect 22252 23364 22256 23420
rect 22192 23360 22256 23364
rect 26952 23420 27016 23424
rect 26952 23364 26956 23420
rect 26956 23364 27012 23420
rect 27012 23364 27016 23420
rect 26952 23360 27016 23364
rect 27032 23420 27096 23424
rect 27032 23364 27036 23420
rect 27036 23364 27092 23420
rect 27092 23364 27096 23420
rect 27032 23360 27096 23364
rect 27112 23420 27176 23424
rect 27112 23364 27116 23420
rect 27116 23364 27172 23420
rect 27172 23364 27176 23420
rect 27112 23360 27176 23364
rect 27192 23420 27256 23424
rect 27192 23364 27196 23420
rect 27196 23364 27252 23420
rect 27252 23364 27256 23420
rect 27192 23360 27256 23364
rect 31952 23420 32016 23424
rect 31952 23364 31956 23420
rect 31956 23364 32012 23420
rect 32012 23364 32016 23420
rect 31952 23360 32016 23364
rect 32032 23420 32096 23424
rect 32032 23364 32036 23420
rect 32036 23364 32092 23420
rect 32092 23364 32096 23420
rect 32032 23360 32096 23364
rect 32112 23420 32176 23424
rect 32112 23364 32116 23420
rect 32116 23364 32172 23420
rect 32172 23364 32176 23420
rect 32112 23360 32176 23364
rect 32192 23420 32256 23424
rect 32192 23364 32196 23420
rect 32196 23364 32252 23420
rect 32252 23364 32256 23420
rect 32192 23360 32256 23364
rect 36952 23420 37016 23424
rect 36952 23364 36956 23420
rect 36956 23364 37012 23420
rect 37012 23364 37016 23420
rect 36952 23360 37016 23364
rect 37032 23420 37096 23424
rect 37032 23364 37036 23420
rect 37036 23364 37092 23420
rect 37092 23364 37096 23420
rect 37032 23360 37096 23364
rect 37112 23420 37176 23424
rect 37112 23364 37116 23420
rect 37116 23364 37172 23420
rect 37172 23364 37176 23420
rect 37112 23360 37176 23364
rect 37192 23420 37256 23424
rect 37192 23364 37196 23420
rect 37196 23364 37252 23420
rect 37252 23364 37256 23420
rect 37192 23360 37256 23364
rect 2612 22876 2676 22880
rect 2612 22820 2616 22876
rect 2616 22820 2672 22876
rect 2672 22820 2676 22876
rect 2612 22816 2676 22820
rect 2692 22876 2756 22880
rect 2692 22820 2696 22876
rect 2696 22820 2752 22876
rect 2752 22820 2756 22876
rect 2692 22816 2756 22820
rect 2772 22876 2836 22880
rect 2772 22820 2776 22876
rect 2776 22820 2832 22876
rect 2832 22820 2836 22876
rect 2772 22816 2836 22820
rect 2852 22876 2916 22880
rect 2852 22820 2856 22876
rect 2856 22820 2912 22876
rect 2912 22820 2916 22876
rect 2852 22816 2916 22820
rect 7612 22876 7676 22880
rect 7612 22820 7616 22876
rect 7616 22820 7672 22876
rect 7672 22820 7676 22876
rect 7612 22816 7676 22820
rect 7692 22876 7756 22880
rect 7692 22820 7696 22876
rect 7696 22820 7752 22876
rect 7752 22820 7756 22876
rect 7692 22816 7756 22820
rect 7772 22876 7836 22880
rect 7772 22820 7776 22876
rect 7776 22820 7832 22876
rect 7832 22820 7836 22876
rect 7772 22816 7836 22820
rect 7852 22876 7916 22880
rect 7852 22820 7856 22876
rect 7856 22820 7912 22876
rect 7912 22820 7916 22876
rect 7852 22816 7916 22820
rect 12612 22876 12676 22880
rect 12612 22820 12616 22876
rect 12616 22820 12672 22876
rect 12672 22820 12676 22876
rect 12612 22816 12676 22820
rect 12692 22876 12756 22880
rect 12692 22820 12696 22876
rect 12696 22820 12752 22876
rect 12752 22820 12756 22876
rect 12692 22816 12756 22820
rect 12772 22876 12836 22880
rect 12772 22820 12776 22876
rect 12776 22820 12832 22876
rect 12832 22820 12836 22876
rect 12772 22816 12836 22820
rect 12852 22876 12916 22880
rect 12852 22820 12856 22876
rect 12856 22820 12912 22876
rect 12912 22820 12916 22876
rect 12852 22816 12916 22820
rect 17612 22876 17676 22880
rect 17612 22820 17616 22876
rect 17616 22820 17672 22876
rect 17672 22820 17676 22876
rect 17612 22816 17676 22820
rect 17692 22876 17756 22880
rect 17692 22820 17696 22876
rect 17696 22820 17752 22876
rect 17752 22820 17756 22876
rect 17692 22816 17756 22820
rect 17772 22876 17836 22880
rect 17772 22820 17776 22876
rect 17776 22820 17832 22876
rect 17832 22820 17836 22876
rect 17772 22816 17836 22820
rect 17852 22876 17916 22880
rect 17852 22820 17856 22876
rect 17856 22820 17912 22876
rect 17912 22820 17916 22876
rect 17852 22816 17916 22820
rect 22612 22876 22676 22880
rect 22612 22820 22616 22876
rect 22616 22820 22672 22876
rect 22672 22820 22676 22876
rect 22612 22816 22676 22820
rect 22692 22876 22756 22880
rect 22692 22820 22696 22876
rect 22696 22820 22752 22876
rect 22752 22820 22756 22876
rect 22692 22816 22756 22820
rect 22772 22876 22836 22880
rect 22772 22820 22776 22876
rect 22776 22820 22832 22876
rect 22832 22820 22836 22876
rect 22772 22816 22836 22820
rect 22852 22876 22916 22880
rect 22852 22820 22856 22876
rect 22856 22820 22912 22876
rect 22912 22820 22916 22876
rect 22852 22816 22916 22820
rect 27612 22876 27676 22880
rect 27612 22820 27616 22876
rect 27616 22820 27672 22876
rect 27672 22820 27676 22876
rect 27612 22816 27676 22820
rect 27692 22876 27756 22880
rect 27692 22820 27696 22876
rect 27696 22820 27752 22876
rect 27752 22820 27756 22876
rect 27692 22816 27756 22820
rect 27772 22876 27836 22880
rect 27772 22820 27776 22876
rect 27776 22820 27832 22876
rect 27832 22820 27836 22876
rect 27772 22816 27836 22820
rect 27852 22876 27916 22880
rect 27852 22820 27856 22876
rect 27856 22820 27912 22876
rect 27912 22820 27916 22876
rect 27852 22816 27916 22820
rect 32612 22876 32676 22880
rect 32612 22820 32616 22876
rect 32616 22820 32672 22876
rect 32672 22820 32676 22876
rect 32612 22816 32676 22820
rect 32692 22876 32756 22880
rect 32692 22820 32696 22876
rect 32696 22820 32752 22876
rect 32752 22820 32756 22876
rect 32692 22816 32756 22820
rect 32772 22876 32836 22880
rect 32772 22820 32776 22876
rect 32776 22820 32832 22876
rect 32832 22820 32836 22876
rect 32772 22816 32836 22820
rect 32852 22876 32916 22880
rect 32852 22820 32856 22876
rect 32856 22820 32912 22876
rect 32912 22820 32916 22876
rect 32852 22816 32916 22820
rect 37612 22876 37676 22880
rect 37612 22820 37616 22876
rect 37616 22820 37672 22876
rect 37672 22820 37676 22876
rect 37612 22816 37676 22820
rect 37692 22876 37756 22880
rect 37692 22820 37696 22876
rect 37696 22820 37752 22876
rect 37752 22820 37756 22876
rect 37692 22816 37756 22820
rect 37772 22876 37836 22880
rect 37772 22820 37776 22876
rect 37776 22820 37832 22876
rect 37832 22820 37836 22876
rect 37772 22816 37836 22820
rect 37852 22876 37916 22880
rect 37852 22820 37856 22876
rect 37856 22820 37912 22876
rect 37912 22820 37916 22876
rect 37852 22816 37916 22820
rect 1952 22332 2016 22336
rect 1952 22276 1956 22332
rect 1956 22276 2012 22332
rect 2012 22276 2016 22332
rect 1952 22272 2016 22276
rect 2032 22332 2096 22336
rect 2032 22276 2036 22332
rect 2036 22276 2092 22332
rect 2092 22276 2096 22332
rect 2032 22272 2096 22276
rect 2112 22332 2176 22336
rect 2112 22276 2116 22332
rect 2116 22276 2172 22332
rect 2172 22276 2176 22332
rect 2112 22272 2176 22276
rect 2192 22332 2256 22336
rect 2192 22276 2196 22332
rect 2196 22276 2252 22332
rect 2252 22276 2256 22332
rect 2192 22272 2256 22276
rect 6952 22332 7016 22336
rect 6952 22276 6956 22332
rect 6956 22276 7012 22332
rect 7012 22276 7016 22332
rect 6952 22272 7016 22276
rect 7032 22332 7096 22336
rect 7032 22276 7036 22332
rect 7036 22276 7092 22332
rect 7092 22276 7096 22332
rect 7032 22272 7096 22276
rect 7112 22332 7176 22336
rect 7112 22276 7116 22332
rect 7116 22276 7172 22332
rect 7172 22276 7176 22332
rect 7112 22272 7176 22276
rect 7192 22332 7256 22336
rect 7192 22276 7196 22332
rect 7196 22276 7252 22332
rect 7252 22276 7256 22332
rect 7192 22272 7256 22276
rect 11952 22332 12016 22336
rect 11952 22276 11956 22332
rect 11956 22276 12012 22332
rect 12012 22276 12016 22332
rect 11952 22272 12016 22276
rect 12032 22332 12096 22336
rect 12032 22276 12036 22332
rect 12036 22276 12092 22332
rect 12092 22276 12096 22332
rect 12032 22272 12096 22276
rect 12112 22332 12176 22336
rect 12112 22276 12116 22332
rect 12116 22276 12172 22332
rect 12172 22276 12176 22332
rect 12112 22272 12176 22276
rect 12192 22332 12256 22336
rect 12192 22276 12196 22332
rect 12196 22276 12252 22332
rect 12252 22276 12256 22332
rect 12192 22272 12256 22276
rect 16952 22332 17016 22336
rect 16952 22276 16956 22332
rect 16956 22276 17012 22332
rect 17012 22276 17016 22332
rect 16952 22272 17016 22276
rect 17032 22332 17096 22336
rect 17032 22276 17036 22332
rect 17036 22276 17092 22332
rect 17092 22276 17096 22332
rect 17032 22272 17096 22276
rect 17112 22332 17176 22336
rect 17112 22276 17116 22332
rect 17116 22276 17172 22332
rect 17172 22276 17176 22332
rect 17112 22272 17176 22276
rect 17192 22332 17256 22336
rect 17192 22276 17196 22332
rect 17196 22276 17252 22332
rect 17252 22276 17256 22332
rect 17192 22272 17256 22276
rect 21952 22332 22016 22336
rect 21952 22276 21956 22332
rect 21956 22276 22012 22332
rect 22012 22276 22016 22332
rect 21952 22272 22016 22276
rect 22032 22332 22096 22336
rect 22032 22276 22036 22332
rect 22036 22276 22092 22332
rect 22092 22276 22096 22332
rect 22032 22272 22096 22276
rect 22112 22332 22176 22336
rect 22112 22276 22116 22332
rect 22116 22276 22172 22332
rect 22172 22276 22176 22332
rect 22112 22272 22176 22276
rect 22192 22332 22256 22336
rect 22192 22276 22196 22332
rect 22196 22276 22252 22332
rect 22252 22276 22256 22332
rect 22192 22272 22256 22276
rect 26952 22332 27016 22336
rect 26952 22276 26956 22332
rect 26956 22276 27012 22332
rect 27012 22276 27016 22332
rect 26952 22272 27016 22276
rect 27032 22332 27096 22336
rect 27032 22276 27036 22332
rect 27036 22276 27092 22332
rect 27092 22276 27096 22332
rect 27032 22272 27096 22276
rect 27112 22332 27176 22336
rect 27112 22276 27116 22332
rect 27116 22276 27172 22332
rect 27172 22276 27176 22332
rect 27112 22272 27176 22276
rect 27192 22332 27256 22336
rect 27192 22276 27196 22332
rect 27196 22276 27252 22332
rect 27252 22276 27256 22332
rect 27192 22272 27256 22276
rect 31952 22332 32016 22336
rect 31952 22276 31956 22332
rect 31956 22276 32012 22332
rect 32012 22276 32016 22332
rect 31952 22272 32016 22276
rect 32032 22332 32096 22336
rect 32032 22276 32036 22332
rect 32036 22276 32092 22332
rect 32092 22276 32096 22332
rect 32032 22272 32096 22276
rect 32112 22332 32176 22336
rect 32112 22276 32116 22332
rect 32116 22276 32172 22332
rect 32172 22276 32176 22332
rect 32112 22272 32176 22276
rect 32192 22332 32256 22336
rect 32192 22276 32196 22332
rect 32196 22276 32252 22332
rect 32252 22276 32256 22332
rect 32192 22272 32256 22276
rect 36952 22332 37016 22336
rect 36952 22276 36956 22332
rect 36956 22276 37012 22332
rect 37012 22276 37016 22332
rect 36952 22272 37016 22276
rect 37032 22332 37096 22336
rect 37032 22276 37036 22332
rect 37036 22276 37092 22332
rect 37092 22276 37096 22332
rect 37032 22272 37096 22276
rect 37112 22332 37176 22336
rect 37112 22276 37116 22332
rect 37116 22276 37172 22332
rect 37172 22276 37176 22332
rect 37112 22272 37176 22276
rect 37192 22332 37256 22336
rect 37192 22276 37196 22332
rect 37196 22276 37252 22332
rect 37252 22276 37256 22332
rect 37192 22272 37256 22276
rect 2612 21788 2676 21792
rect 2612 21732 2616 21788
rect 2616 21732 2672 21788
rect 2672 21732 2676 21788
rect 2612 21728 2676 21732
rect 2692 21788 2756 21792
rect 2692 21732 2696 21788
rect 2696 21732 2752 21788
rect 2752 21732 2756 21788
rect 2692 21728 2756 21732
rect 2772 21788 2836 21792
rect 2772 21732 2776 21788
rect 2776 21732 2832 21788
rect 2832 21732 2836 21788
rect 2772 21728 2836 21732
rect 2852 21788 2916 21792
rect 2852 21732 2856 21788
rect 2856 21732 2912 21788
rect 2912 21732 2916 21788
rect 2852 21728 2916 21732
rect 7612 21788 7676 21792
rect 7612 21732 7616 21788
rect 7616 21732 7672 21788
rect 7672 21732 7676 21788
rect 7612 21728 7676 21732
rect 7692 21788 7756 21792
rect 7692 21732 7696 21788
rect 7696 21732 7752 21788
rect 7752 21732 7756 21788
rect 7692 21728 7756 21732
rect 7772 21788 7836 21792
rect 7772 21732 7776 21788
rect 7776 21732 7832 21788
rect 7832 21732 7836 21788
rect 7772 21728 7836 21732
rect 7852 21788 7916 21792
rect 7852 21732 7856 21788
rect 7856 21732 7912 21788
rect 7912 21732 7916 21788
rect 7852 21728 7916 21732
rect 12612 21788 12676 21792
rect 12612 21732 12616 21788
rect 12616 21732 12672 21788
rect 12672 21732 12676 21788
rect 12612 21728 12676 21732
rect 12692 21788 12756 21792
rect 12692 21732 12696 21788
rect 12696 21732 12752 21788
rect 12752 21732 12756 21788
rect 12692 21728 12756 21732
rect 12772 21788 12836 21792
rect 12772 21732 12776 21788
rect 12776 21732 12832 21788
rect 12832 21732 12836 21788
rect 12772 21728 12836 21732
rect 12852 21788 12916 21792
rect 12852 21732 12856 21788
rect 12856 21732 12912 21788
rect 12912 21732 12916 21788
rect 12852 21728 12916 21732
rect 17612 21788 17676 21792
rect 17612 21732 17616 21788
rect 17616 21732 17672 21788
rect 17672 21732 17676 21788
rect 17612 21728 17676 21732
rect 17692 21788 17756 21792
rect 17692 21732 17696 21788
rect 17696 21732 17752 21788
rect 17752 21732 17756 21788
rect 17692 21728 17756 21732
rect 17772 21788 17836 21792
rect 17772 21732 17776 21788
rect 17776 21732 17832 21788
rect 17832 21732 17836 21788
rect 17772 21728 17836 21732
rect 17852 21788 17916 21792
rect 17852 21732 17856 21788
rect 17856 21732 17912 21788
rect 17912 21732 17916 21788
rect 17852 21728 17916 21732
rect 22612 21788 22676 21792
rect 22612 21732 22616 21788
rect 22616 21732 22672 21788
rect 22672 21732 22676 21788
rect 22612 21728 22676 21732
rect 22692 21788 22756 21792
rect 22692 21732 22696 21788
rect 22696 21732 22752 21788
rect 22752 21732 22756 21788
rect 22692 21728 22756 21732
rect 22772 21788 22836 21792
rect 22772 21732 22776 21788
rect 22776 21732 22832 21788
rect 22832 21732 22836 21788
rect 22772 21728 22836 21732
rect 22852 21788 22916 21792
rect 22852 21732 22856 21788
rect 22856 21732 22912 21788
rect 22912 21732 22916 21788
rect 22852 21728 22916 21732
rect 27612 21788 27676 21792
rect 27612 21732 27616 21788
rect 27616 21732 27672 21788
rect 27672 21732 27676 21788
rect 27612 21728 27676 21732
rect 27692 21788 27756 21792
rect 27692 21732 27696 21788
rect 27696 21732 27752 21788
rect 27752 21732 27756 21788
rect 27692 21728 27756 21732
rect 27772 21788 27836 21792
rect 27772 21732 27776 21788
rect 27776 21732 27832 21788
rect 27832 21732 27836 21788
rect 27772 21728 27836 21732
rect 27852 21788 27916 21792
rect 27852 21732 27856 21788
rect 27856 21732 27912 21788
rect 27912 21732 27916 21788
rect 27852 21728 27916 21732
rect 32612 21788 32676 21792
rect 32612 21732 32616 21788
rect 32616 21732 32672 21788
rect 32672 21732 32676 21788
rect 32612 21728 32676 21732
rect 32692 21788 32756 21792
rect 32692 21732 32696 21788
rect 32696 21732 32752 21788
rect 32752 21732 32756 21788
rect 32692 21728 32756 21732
rect 32772 21788 32836 21792
rect 32772 21732 32776 21788
rect 32776 21732 32832 21788
rect 32832 21732 32836 21788
rect 32772 21728 32836 21732
rect 32852 21788 32916 21792
rect 32852 21732 32856 21788
rect 32856 21732 32912 21788
rect 32912 21732 32916 21788
rect 32852 21728 32916 21732
rect 37612 21788 37676 21792
rect 37612 21732 37616 21788
rect 37616 21732 37672 21788
rect 37672 21732 37676 21788
rect 37612 21728 37676 21732
rect 37692 21788 37756 21792
rect 37692 21732 37696 21788
rect 37696 21732 37752 21788
rect 37752 21732 37756 21788
rect 37692 21728 37756 21732
rect 37772 21788 37836 21792
rect 37772 21732 37776 21788
rect 37776 21732 37832 21788
rect 37832 21732 37836 21788
rect 37772 21728 37836 21732
rect 37852 21788 37916 21792
rect 37852 21732 37856 21788
rect 37856 21732 37912 21788
rect 37912 21732 37916 21788
rect 37852 21728 37916 21732
rect 1952 21244 2016 21248
rect 1952 21188 1956 21244
rect 1956 21188 2012 21244
rect 2012 21188 2016 21244
rect 1952 21184 2016 21188
rect 2032 21244 2096 21248
rect 2032 21188 2036 21244
rect 2036 21188 2092 21244
rect 2092 21188 2096 21244
rect 2032 21184 2096 21188
rect 2112 21244 2176 21248
rect 2112 21188 2116 21244
rect 2116 21188 2172 21244
rect 2172 21188 2176 21244
rect 2112 21184 2176 21188
rect 2192 21244 2256 21248
rect 2192 21188 2196 21244
rect 2196 21188 2252 21244
rect 2252 21188 2256 21244
rect 2192 21184 2256 21188
rect 6952 21244 7016 21248
rect 6952 21188 6956 21244
rect 6956 21188 7012 21244
rect 7012 21188 7016 21244
rect 6952 21184 7016 21188
rect 7032 21244 7096 21248
rect 7032 21188 7036 21244
rect 7036 21188 7092 21244
rect 7092 21188 7096 21244
rect 7032 21184 7096 21188
rect 7112 21244 7176 21248
rect 7112 21188 7116 21244
rect 7116 21188 7172 21244
rect 7172 21188 7176 21244
rect 7112 21184 7176 21188
rect 7192 21244 7256 21248
rect 7192 21188 7196 21244
rect 7196 21188 7252 21244
rect 7252 21188 7256 21244
rect 7192 21184 7256 21188
rect 11952 21244 12016 21248
rect 11952 21188 11956 21244
rect 11956 21188 12012 21244
rect 12012 21188 12016 21244
rect 11952 21184 12016 21188
rect 12032 21244 12096 21248
rect 12032 21188 12036 21244
rect 12036 21188 12092 21244
rect 12092 21188 12096 21244
rect 12032 21184 12096 21188
rect 12112 21244 12176 21248
rect 12112 21188 12116 21244
rect 12116 21188 12172 21244
rect 12172 21188 12176 21244
rect 12112 21184 12176 21188
rect 12192 21244 12256 21248
rect 12192 21188 12196 21244
rect 12196 21188 12252 21244
rect 12252 21188 12256 21244
rect 12192 21184 12256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 21952 21244 22016 21248
rect 21952 21188 21956 21244
rect 21956 21188 22012 21244
rect 22012 21188 22016 21244
rect 21952 21184 22016 21188
rect 22032 21244 22096 21248
rect 22032 21188 22036 21244
rect 22036 21188 22092 21244
rect 22092 21188 22096 21244
rect 22032 21184 22096 21188
rect 22112 21244 22176 21248
rect 22112 21188 22116 21244
rect 22116 21188 22172 21244
rect 22172 21188 22176 21244
rect 22112 21184 22176 21188
rect 22192 21244 22256 21248
rect 22192 21188 22196 21244
rect 22196 21188 22252 21244
rect 22252 21188 22256 21244
rect 22192 21184 22256 21188
rect 26952 21244 27016 21248
rect 26952 21188 26956 21244
rect 26956 21188 27012 21244
rect 27012 21188 27016 21244
rect 26952 21184 27016 21188
rect 27032 21244 27096 21248
rect 27032 21188 27036 21244
rect 27036 21188 27092 21244
rect 27092 21188 27096 21244
rect 27032 21184 27096 21188
rect 27112 21244 27176 21248
rect 27112 21188 27116 21244
rect 27116 21188 27172 21244
rect 27172 21188 27176 21244
rect 27112 21184 27176 21188
rect 27192 21244 27256 21248
rect 27192 21188 27196 21244
rect 27196 21188 27252 21244
rect 27252 21188 27256 21244
rect 27192 21184 27256 21188
rect 31952 21244 32016 21248
rect 31952 21188 31956 21244
rect 31956 21188 32012 21244
rect 32012 21188 32016 21244
rect 31952 21184 32016 21188
rect 32032 21244 32096 21248
rect 32032 21188 32036 21244
rect 32036 21188 32092 21244
rect 32092 21188 32096 21244
rect 32032 21184 32096 21188
rect 32112 21244 32176 21248
rect 32112 21188 32116 21244
rect 32116 21188 32172 21244
rect 32172 21188 32176 21244
rect 32112 21184 32176 21188
rect 32192 21244 32256 21248
rect 32192 21188 32196 21244
rect 32196 21188 32252 21244
rect 32252 21188 32256 21244
rect 32192 21184 32256 21188
rect 36952 21244 37016 21248
rect 36952 21188 36956 21244
rect 36956 21188 37012 21244
rect 37012 21188 37016 21244
rect 36952 21184 37016 21188
rect 37032 21244 37096 21248
rect 37032 21188 37036 21244
rect 37036 21188 37092 21244
rect 37092 21188 37096 21244
rect 37032 21184 37096 21188
rect 37112 21244 37176 21248
rect 37112 21188 37116 21244
rect 37116 21188 37172 21244
rect 37172 21188 37176 21244
rect 37112 21184 37176 21188
rect 37192 21244 37256 21248
rect 37192 21188 37196 21244
rect 37196 21188 37252 21244
rect 37252 21188 37256 21244
rect 37192 21184 37256 21188
rect 2612 20700 2676 20704
rect 2612 20644 2616 20700
rect 2616 20644 2672 20700
rect 2672 20644 2676 20700
rect 2612 20640 2676 20644
rect 2692 20700 2756 20704
rect 2692 20644 2696 20700
rect 2696 20644 2752 20700
rect 2752 20644 2756 20700
rect 2692 20640 2756 20644
rect 2772 20700 2836 20704
rect 2772 20644 2776 20700
rect 2776 20644 2832 20700
rect 2832 20644 2836 20700
rect 2772 20640 2836 20644
rect 2852 20700 2916 20704
rect 2852 20644 2856 20700
rect 2856 20644 2912 20700
rect 2912 20644 2916 20700
rect 2852 20640 2916 20644
rect 7612 20700 7676 20704
rect 7612 20644 7616 20700
rect 7616 20644 7672 20700
rect 7672 20644 7676 20700
rect 7612 20640 7676 20644
rect 7692 20700 7756 20704
rect 7692 20644 7696 20700
rect 7696 20644 7752 20700
rect 7752 20644 7756 20700
rect 7692 20640 7756 20644
rect 7772 20700 7836 20704
rect 7772 20644 7776 20700
rect 7776 20644 7832 20700
rect 7832 20644 7836 20700
rect 7772 20640 7836 20644
rect 7852 20700 7916 20704
rect 7852 20644 7856 20700
rect 7856 20644 7912 20700
rect 7912 20644 7916 20700
rect 7852 20640 7916 20644
rect 12612 20700 12676 20704
rect 12612 20644 12616 20700
rect 12616 20644 12672 20700
rect 12672 20644 12676 20700
rect 12612 20640 12676 20644
rect 12692 20700 12756 20704
rect 12692 20644 12696 20700
rect 12696 20644 12752 20700
rect 12752 20644 12756 20700
rect 12692 20640 12756 20644
rect 12772 20700 12836 20704
rect 12772 20644 12776 20700
rect 12776 20644 12832 20700
rect 12832 20644 12836 20700
rect 12772 20640 12836 20644
rect 12852 20700 12916 20704
rect 12852 20644 12856 20700
rect 12856 20644 12912 20700
rect 12912 20644 12916 20700
rect 12852 20640 12916 20644
rect 17612 20700 17676 20704
rect 17612 20644 17616 20700
rect 17616 20644 17672 20700
rect 17672 20644 17676 20700
rect 17612 20640 17676 20644
rect 17692 20700 17756 20704
rect 17692 20644 17696 20700
rect 17696 20644 17752 20700
rect 17752 20644 17756 20700
rect 17692 20640 17756 20644
rect 17772 20700 17836 20704
rect 17772 20644 17776 20700
rect 17776 20644 17832 20700
rect 17832 20644 17836 20700
rect 17772 20640 17836 20644
rect 17852 20700 17916 20704
rect 17852 20644 17856 20700
rect 17856 20644 17912 20700
rect 17912 20644 17916 20700
rect 17852 20640 17916 20644
rect 22612 20700 22676 20704
rect 22612 20644 22616 20700
rect 22616 20644 22672 20700
rect 22672 20644 22676 20700
rect 22612 20640 22676 20644
rect 22692 20700 22756 20704
rect 22692 20644 22696 20700
rect 22696 20644 22752 20700
rect 22752 20644 22756 20700
rect 22692 20640 22756 20644
rect 22772 20700 22836 20704
rect 22772 20644 22776 20700
rect 22776 20644 22832 20700
rect 22832 20644 22836 20700
rect 22772 20640 22836 20644
rect 22852 20700 22916 20704
rect 22852 20644 22856 20700
rect 22856 20644 22912 20700
rect 22912 20644 22916 20700
rect 22852 20640 22916 20644
rect 27612 20700 27676 20704
rect 27612 20644 27616 20700
rect 27616 20644 27672 20700
rect 27672 20644 27676 20700
rect 27612 20640 27676 20644
rect 27692 20700 27756 20704
rect 27692 20644 27696 20700
rect 27696 20644 27752 20700
rect 27752 20644 27756 20700
rect 27692 20640 27756 20644
rect 27772 20700 27836 20704
rect 27772 20644 27776 20700
rect 27776 20644 27832 20700
rect 27832 20644 27836 20700
rect 27772 20640 27836 20644
rect 27852 20700 27916 20704
rect 27852 20644 27856 20700
rect 27856 20644 27912 20700
rect 27912 20644 27916 20700
rect 27852 20640 27916 20644
rect 32612 20700 32676 20704
rect 32612 20644 32616 20700
rect 32616 20644 32672 20700
rect 32672 20644 32676 20700
rect 32612 20640 32676 20644
rect 32692 20700 32756 20704
rect 32692 20644 32696 20700
rect 32696 20644 32752 20700
rect 32752 20644 32756 20700
rect 32692 20640 32756 20644
rect 32772 20700 32836 20704
rect 32772 20644 32776 20700
rect 32776 20644 32832 20700
rect 32832 20644 32836 20700
rect 32772 20640 32836 20644
rect 32852 20700 32916 20704
rect 32852 20644 32856 20700
rect 32856 20644 32912 20700
rect 32912 20644 32916 20700
rect 32852 20640 32916 20644
rect 37612 20700 37676 20704
rect 37612 20644 37616 20700
rect 37616 20644 37672 20700
rect 37672 20644 37676 20700
rect 37612 20640 37676 20644
rect 37692 20700 37756 20704
rect 37692 20644 37696 20700
rect 37696 20644 37752 20700
rect 37752 20644 37756 20700
rect 37692 20640 37756 20644
rect 37772 20700 37836 20704
rect 37772 20644 37776 20700
rect 37776 20644 37832 20700
rect 37832 20644 37836 20700
rect 37772 20640 37836 20644
rect 37852 20700 37916 20704
rect 37852 20644 37856 20700
rect 37856 20644 37912 20700
rect 37912 20644 37916 20700
rect 37852 20640 37916 20644
rect 1952 20156 2016 20160
rect 1952 20100 1956 20156
rect 1956 20100 2012 20156
rect 2012 20100 2016 20156
rect 1952 20096 2016 20100
rect 2032 20156 2096 20160
rect 2032 20100 2036 20156
rect 2036 20100 2092 20156
rect 2092 20100 2096 20156
rect 2032 20096 2096 20100
rect 2112 20156 2176 20160
rect 2112 20100 2116 20156
rect 2116 20100 2172 20156
rect 2172 20100 2176 20156
rect 2112 20096 2176 20100
rect 2192 20156 2256 20160
rect 2192 20100 2196 20156
rect 2196 20100 2252 20156
rect 2252 20100 2256 20156
rect 2192 20096 2256 20100
rect 6952 20156 7016 20160
rect 6952 20100 6956 20156
rect 6956 20100 7012 20156
rect 7012 20100 7016 20156
rect 6952 20096 7016 20100
rect 7032 20156 7096 20160
rect 7032 20100 7036 20156
rect 7036 20100 7092 20156
rect 7092 20100 7096 20156
rect 7032 20096 7096 20100
rect 7112 20156 7176 20160
rect 7112 20100 7116 20156
rect 7116 20100 7172 20156
rect 7172 20100 7176 20156
rect 7112 20096 7176 20100
rect 7192 20156 7256 20160
rect 7192 20100 7196 20156
rect 7196 20100 7252 20156
rect 7252 20100 7256 20156
rect 7192 20096 7256 20100
rect 11952 20156 12016 20160
rect 11952 20100 11956 20156
rect 11956 20100 12012 20156
rect 12012 20100 12016 20156
rect 11952 20096 12016 20100
rect 12032 20156 12096 20160
rect 12032 20100 12036 20156
rect 12036 20100 12092 20156
rect 12092 20100 12096 20156
rect 12032 20096 12096 20100
rect 12112 20156 12176 20160
rect 12112 20100 12116 20156
rect 12116 20100 12172 20156
rect 12172 20100 12176 20156
rect 12112 20096 12176 20100
rect 12192 20156 12256 20160
rect 12192 20100 12196 20156
rect 12196 20100 12252 20156
rect 12252 20100 12256 20156
rect 12192 20096 12256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 21952 20156 22016 20160
rect 21952 20100 21956 20156
rect 21956 20100 22012 20156
rect 22012 20100 22016 20156
rect 21952 20096 22016 20100
rect 22032 20156 22096 20160
rect 22032 20100 22036 20156
rect 22036 20100 22092 20156
rect 22092 20100 22096 20156
rect 22032 20096 22096 20100
rect 22112 20156 22176 20160
rect 22112 20100 22116 20156
rect 22116 20100 22172 20156
rect 22172 20100 22176 20156
rect 22112 20096 22176 20100
rect 22192 20156 22256 20160
rect 22192 20100 22196 20156
rect 22196 20100 22252 20156
rect 22252 20100 22256 20156
rect 22192 20096 22256 20100
rect 26952 20156 27016 20160
rect 26952 20100 26956 20156
rect 26956 20100 27012 20156
rect 27012 20100 27016 20156
rect 26952 20096 27016 20100
rect 27032 20156 27096 20160
rect 27032 20100 27036 20156
rect 27036 20100 27092 20156
rect 27092 20100 27096 20156
rect 27032 20096 27096 20100
rect 27112 20156 27176 20160
rect 27112 20100 27116 20156
rect 27116 20100 27172 20156
rect 27172 20100 27176 20156
rect 27112 20096 27176 20100
rect 27192 20156 27256 20160
rect 27192 20100 27196 20156
rect 27196 20100 27252 20156
rect 27252 20100 27256 20156
rect 27192 20096 27256 20100
rect 31952 20156 32016 20160
rect 31952 20100 31956 20156
rect 31956 20100 32012 20156
rect 32012 20100 32016 20156
rect 31952 20096 32016 20100
rect 32032 20156 32096 20160
rect 32032 20100 32036 20156
rect 32036 20100 32092 20156
rect 32092 20100 32096 20156
rect 32032 20096 32096 20100
rect 32112 20156 32176 20160
rect 32112 20100 32116 20156
rect 32116 20100 32172 20156
rect 32172 20100 32176 20156
rect 32112 20096 32176 20100
rect 32192 20156 32256 20160
rect 32192 20100 32196 20156
rect 32196 20100 32252 20156
rect 32252 20100 32256 20156
rect 32192 20096 32256 20100
rect 36952 20156 37016 20160
rect 36952 20100 36956 20156
rect 36956 20100 37012 20156
rect 37012 20100 37016 20156
rect 36952 20096 37016 20100
rect 37032 20156 37096 20160
rect 37032 20100 37036 20156
rect 37036 20100 37092 20156
rect 37092 20100 37096 20156
rect 37032 20096 37096 20100
rect 37112 20156 37176 20160
rect 37112 20100 37116 20156
rect 37116 20100 37172 20156
rect 37172 20100 37176 20156
rect 37112 20096 37176 20100
rect 37192 20156 37256 20160
rect 37192 20100 37196 20156
rect 37196 20100 37252 20156
rect 37252 20100 37256 20156
rect 37192 20096 37256 20100
rect 2612 19612 2676 19616
rect 2612 19556 2616 19612
rect 2616 19556 2672 19612
rect 2672 19556 2676 19612
rect 2612 19552 2676 19556
rect 2692 19612 2756 19616
rect 2692 19556 2696 19612
rect 2696 19556 2752 19612
rect 2752 19556 2756 19612
rect 2692 19552 2756 19556
rect 2772 19612 2836 19616
rect 2772 19556 2776 19612
rect 2776 19556 2832 19612
rect 2832 19556 2836 19612
rect 2772 19552 2836 19556
rect 2852 19612 2916 19616
rect 2852 19556 2856 19612
rect 2856 19556 2912 19612
rect 2912 19556 2916 19612
rect 2852 19552 2916 19556
rect 7612 19612 7676 19616
rect 7612 19556 7616 19612
rect 7616 19556 7672 19612
rect 7672 19556 7676 19612
rect 7612 19552 7676 19556
rect 7692 19612 7756 19616
rect 7692 19556 7696 19612
rect 7696 19556 7752 19612
rect 7752 19556 7756 19612
rect 7692 19552 7756 19556
rect 7772 19612 7836 19616
rect 7772 19556 7776 19612
rect 7776 19556 7832 19612
rect 7832 19556 7836 19612
rect 7772 19552 7836 19556
rect 7852 19612 7916 19616
rect 7852 19556 7856 19612
rect 7856 19556 7912 19612
rect 7912 19556 7916 19612
rect 7852 19552 7916 19556
rect 12612 19612 12676 19616
rect 12612 19556 12616 19612
rect 12616 19556 12672 19612
rect 12672 19556 12676 19612
rect 12612 19552 12676 19556
rect 12692 19612 12756 19616
rect 12692 19556 12696 19612
rect 12696 19556 12752 19612
rect 12752 19556 12756 19612
rect 12692 19552 12756 19556
rect 12772 19612 12836 19616
rect 12772 19556 12776 19612
rect 12776 19556 12832 19612
rect 12832 19556 12836 19612
rect 12772 19552 12836 19556
rect 12852 19612 12916 19616
rect 12852 19556 12856 19612
rect 12856 19556 12912 19612
rect 12912 19556 12916 19612
rect 12852 19552 12916 19556
rect 17612 19612 17676 19616
rect 17612 19556 17616 19612
rect 17616 19556 17672 19612
rect 17672 19556 17676 19612
rect 17612 19552 17676 19556
rect 17692 19612 17756 19616
rect 17692 19556 17696 19612
rect 17696 19556 17752 19612
rect 17752 19556 17756 19612
rect 17692 19552 17756 19556
rect 17772 19612 17836 19616
rect 17772 19556 17776 19612
rect 17776 19556 17832 19612
rect 17832 19556 17836 19612
rect 17772 19552 17836 19556
rect 17852 19612 17916 19616
rect 17852 19556 17856 19612
rect 17856 19556 17912 19612
rect 17912 19556 17916 19612
rect 17852 19552 17916 19556
rect 22612 19612 22676 19616
rect 22612 19556 22616 19612
rect 22616 19556 22672 19612
rect 22672 19556 22676 19612
rect 22612 19552 22676 19556
rect 22692 19612 22756 19616
rect 22692 19556 22696 19612
rect 22696 19556 22752 19612
rect 22752 19556 22756 19612
rect 22692 19552 22756 19556
rect 22772 19612 22836 19616
rect 22772 19556 22776 19612
rect 22776 19556 22832 19612
rect 22832 19556 22836 19612
rect 22772 19552 22836 19556
rect 22852 19612 22916 19616
rect 22852 19556 22856 19612
rect 22856 19556 22912 19612
rect 22912 19556 22916 19612
rect 22852 19552 22916 19556
rect 27612 19612 27676 19616
rect 27612 19556 27616 19612
rect 27616 19556 27672 19612
rect 27672 19556 27676 19612
rect 27612 19552 27676 19556
rect 27692 19612 27756 19616
rect 27692 19556 27696 19612
rect 27696 19556 27752 19612
rect 27752 19556 27756 19612
rect 27692 19552 27756 19556
rect 27772 19612 27836 19616
rect 27772 19556 27776 19612
rect 27776 19556 27832 19612
rect 27832 19556 27836 19612
rect 27772 19552 27836 19556
rect 27852 19612 27916 19616
rect 27852 19556 27856 19612
rect 27856 19556 27912 19612
rect 27912 19556 27916 19612
rect 27852 19552 27916 19556
rect 32612 19612 32676 19616
rect 32612 19556 32616 19612
rect 32616 19556 32672 19612
rect 32672 19556 32676 19612
rect 32612 19552 32676 19556
rect 32692 19612 32756 19616
rect 32692 19556 32696 19612
rect 32696 19556 32752 19612
rect 32752 19556 32756 19612
rect 32692 19552 32756 19556
rect 32772 19612 32836 19616
rect 32772 19556 32776 19612
rect 32776 19556 32832 19612
rect 32832 19556 32836 19612
rect 32772 19552 32836 19556
rect 32852 19612 32916 19616
rect 32852 19556 32856 19612
rect 32856 19556 32912 19612
rect 32912 19556 32916 19612
rect 32852 19552 32916 19556
rect 37612 19612 37676 19616
rect 37612 19556 37616 19612
rect 37616 19556 37672 19612
rect 37672 19556 37676 19612
rect 37612 19552 37676 19556
rect 37692 19612 37756 19616
rect 37692 19556 37696 19612
rect 37696 19556 37752 19612
rect 37752 19556 37756 19612
rect 37692 19552 37756 19556
rect 37772 19612 37836 19616
rect 37772 19556 37776 19612
rect 37776 19556 37832 19612
rect 37832 19556 37836 19612
rect 37772 19552 37836 19556
rect 37852 19612 37916 19616
rect 37852 19556 37856 19612
rect 37856 19556 37912 19612
rect 37912 19556 37916 19612
rect 37852 19552 37916 19556
rect 1952 19068 2016 19072
rect 1952 19012 1956 19068
rect 1956 19012 2012 19068
rect 2012 19012 2016 19068
rect 1952 19008 2016 19012
rect 2032 19068 2096 19072
rect 2032 19012 2036 19068
rect 2036 19012 2092 19068
rect 2092 19012 2096 19068
rect 2032 19008 2096 19012
rect 2112 19068 2176 19072
rect 2112 19012 2116 19068
rect 2116 19012 2172 19068
rect 2172 19012 2176 19068
rect 2112 19008 2176 19012
rect 2192 19068 2256 19072
rect 2192 19012 2196 19068
rect 2196 19012 2252 19068
rect 2252 19012 2256 19068
rect 2192 19008 2256 19012
rect 6952 19068 7016 19072
rect 6952 19012 6956 19068
rect 6956 19012 7012 19068
rect 7012 19012 7016 19068
rect 6952 19008 7016 19012
rect 7032 19068 7096 19072
rect 7032 19012 7036 19068
rect 7036 19012 7092 19068
rect 7092 19012 7096 19068
rect 7032 19008 7096 19012
rect 7112 19068 7176 19072
rect 7112 19012 7116 19068
rect 7116 19012 7172 19068
rect 7172 19012 7176 19068
rect 7112 19008 7176 19012
rect 7192 19068 7256 19072
rect 7192 19012 7196 19068
rect 7196 19012 7252 19068
rect 7252 19012 7256 19068
rect 7192 19008 7256 19012
rect 11952 19068 12016 19072
rect 11952 19012 11956 19068
rect 11956 19012 12012 19068
rect 12012 19012 12016 19068
rect 11952 19008 12016 19012
rect 12032 19068 12096 19072
rect 12032 19012 12036 19068
rect 12036 19012 12092 19068
rect 12092 19012 12096 19068
rect 12032 19008 12096 19012
rect 12112 19068 12176 19072
rect 12112 19012 12116 19068
rect 12116 19012 12172 19068
rect 12172 19012 12176 19068
rect 12112 19008 12176 19012
rect 12192 19068 12256 19072
rect 12192 19012 12196 19068
rect 12196 19012 12252 19068
rect 12252 19012 12256 19068
rect 12192 19008 12256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 21952 19068 22016 19072
rect 21952 19012 21956 19068
rect 21956 19012 22012 19068
rect 22012 19012 22016 19068
rect 21952 19008 22016 19012
rect 22032 19068 22096 19072
rect 22032 19012 22036 19068
rect 22036 19012 22092 19068
rect 22092 19012 22096 19068
rect 22032 19008 22096 19012
rect 22112 19068 22176 19072
rect 22112 19012 22116 19068
rect 22116 19012 22172 19068
rect 22172 19012 22176 19068
rect 22112 19008 22176 19012
rect 22192 19068 22256 19072
rect 22192 19012 22196 19068
rect 22196 19012 22252 19068
rect 22252 19012 22256 19068
rect 22192 19008 22256 19012
rect 26952 19068 27016 19072
rect 26952 19012 26956 19068
rect 26956 19012 27012 19068
rect 27012 19012 27016 19068
rect 26952 19008 27016 19012
rect 27032 19068 27096 19072
rect 27032 19012 27036 19068
rect 27036 19012 27092 19068
rect 27092 19012 27096 19068
rect 27032 19008 27096 19012
rect 27112 19068 27176 19072
rect 27112 19012 27116 19068
rect 27116 19012 27172 19068
rect 27172 19012 27176 19068
rect 27112 19008 27176 19012
rect 27192 19068 27256 19072
rect 27192 19012 27196 19068
rect 27196 19012 27252 19068
rect 27252 19012 27256 19068
rect 27192 19008 27256 19012
rect 31952 19068 32016 19072
rect 31952 19012 31956 19068
rect 31956 19012 32012 19068
rect 32012 19012 32016 19068
rect 31952 19008 32016 19012
rect 32032 19068 32096 19072
rect 32032 19012 32036 19068
rect 32036 19012 32092 19068
rect 32092 19012 32096 19068
rect 32032 19008 32096 19012
rect 32112 19068 32176 19072
rect 32112 19012 32116 19068
rect 32116 19012 32172 19068
rect 32172 19012 32176 19068
rect 32112 19008 32176 19012
rect 32192 19068 32256 19072
rect 32192 19012 32196 19068
rect 32196 19012 32252 19068
rect 32252 19012 32256 19068
rect 32192 19008 32256 19012
rect 36952 19068 37016 19072
rect 36952 19012 36956 19068
rect 36956 19012 37012 19068
rect 37012 19012 37016 19068
rect 36952 19008 37016 19012
rect 37032 19068 37096 19072
rect 37032 19012 37036 19068
rect 37036 19012 37092 19068
rect 37092 19012 37096 19068
rect 37032 19008 37096 19012
rect 37112 19068 37176 19072
rect 37112 19012 37116 19068
rect 37116 19012 37172 19068
rect 37172 19012 37176 19068
rect 37112 19008 37176 19012
rect 37192 19068 37256 19072
rect 37192 19012 37196 19068
rect 37196 19012 37252 19068
rect 37252 19012 37256 19068
rect 37192 19008 37256 19012
rect 2612 18524 2676 18528
rect 2612 18468 2616 18524
rect 2616 18468 2672 18524
rect 2672 18468 2676 18524
rect 2612 18464 2676 18468
rect 2692 18524 2756 18528
rect 2692 18468 2696 18524
rect 2696 18468 2752 18524
rect 2752 18468 2756 18524
rect 2692 18464 2756 18468
rect 2772 18524 2836 18528
rect 2772 18468 2776 18524
rect 2776 18468 2832 18524
rect 2832 18468 2836 18524
rect 2772 18464 2836 18468
rect 2852 18524 2916 18528
rect 2852 18468 2856 18524
rect 2856 18468 2912 18524
rect 2912 18468 2916 18524
rect 2852 18464 2916 18468
rect 7612 18524 7676 18528
rect 7612 18468 7616 18524
rect 7616 18468 7672 18524
rect 7672 18468 7676 18524
rect 7612 18464 7676 18468
rect 7692 18524 7756 18528
rect 7692 18468 7696 18524
rect 7696 18468 7752 18524
rect 7752 18468 7756 18524
rect 7692 18464 7756 18468
rect 7772 18524 7836 18528
rect 7772 18468 7776 18524
rect 7776 18468 7832 18524
rect 7832 18468 7836 18524
rect 7772 18464 7836 18468
rect 7852 18524 7916 18528
rect 7852 18468 7856 18524
rect 7856 18468 7912 18524
rect 7912 18468 7916 18524
rect 7852 18464 7916 18468
rect 12612 18524 12676 18528
rect 12612 18468 12616 18524
rect 12616 18468 12672 18524
rect 12672 18468 12676 18524
rect 12612 18464 12676 18468
rect 12692 18524 12756 18528
rect 12692 18468 12696 18524
rect 12696 18468 12752 18524
rect 12752 18468 12756 18524
rect 12692 18464 12756 18468
rect 12772 18524 12836 18528
rect 12772 18468 12776 18524
rect 12776 18468 12832 18524
rect 12832 18468 12836 18524
rect 12772 18464 12836 18468
rect 12852 18524 12916 18528
rect 12852 18468 12856 18524
rect 12856 18468 12912 18524
rect 12912 18468 12916 18524
rect 12852 18464 12916 18468
rect 17612 18524 17676 18528
rect 17612 18468 17616 18524
rect 17616 18468 17672 18524
rect 17672 18468 17676 18524
rect 17612 18464 17676 18468
rect 17692 18524 17756 18528
rect 17692 18468 17696 18524
rect 17696 18468 17752 18524
rect 17752 18468 17756 18524
rect 17692 18464 17756 18468
rect 17772 18524 17836 18528
rect 17772 18468 17776 18524
rect 17776 18468 17832 18524
rect 17832 18468 17836 18524
rect 17772 18464 17836 18468
rect 17852 18524 17916 18528
rect 17852 18468 17856 18524
rect 17856 18468 17912 18524
rect 17912 18468 17916 18524
rect 17852 18464 17916 18468
rect 22612 18524 22676 18528
rect 22612 18468 22616 18524
rect 22616 18468 22672 18524
rect 22672 18468 22676 18524
rect 22612 18464 22676 18468
rect 22692 18524 22756 18528
rect 22692 18468 22696 18524
rect 22696 18468 22752 18524
rect 22752 18468 22756 18524
rect 22692 18464 22756 18468
rect 22772 18524 22836 18528
rect 22772 18468 22776 18524
rect 22776 18468 22832 18524
rect 22832 18468 22836 18524
rect 22772 18464 22836 18468
rect 22852 18524 22916 18528
rect 22852 18468 22856 18524
rect 22856 18468 22912 18524
rect 22912 18468 22916 18524
rect 22852 18464 22916 18468
rect 27612 18524 27676 18528
rect 27612 18468 27616 18524
rect 27616 18468 27672 18524
rect 27672 18468 27676 18524
rect 27612 18464 27676 18468
rect 27692 18524 27756 18528
rect 27692 18468 27696 18524
rect 27696 18468 27752 18524
rect 27752 18468 27756 18524
rect 27692 18464 27756 18468
rect 27772 18524 27836 18528
rect 27772 18468 27776 18524
rect 27776 18468 27832 18524
rect 27832 18468 27836 18524
rect 27772 18464 27836 18468
rect 27852 18524 27916 18528
rect 27852 18468 27856 18524
rect 27856 18468 27912 18524
rect 27912 18468 27916 18524
rect 27852 18464 27916 18468
rect 32612 18524 32676 18528
rect 32612 18468 32616 18524
rect 32616 18468 32672 18524
rect 32672 18468 32676 18524
rect 32612 18464 32676 18468
rect 32692 18524 32756 18528
rect 32692 18468 32696 18524
rect 32696 18468 32752 18524
rect 32752 18468 32756 18524
rect 32692 18464 32756 18468
rect 32772 18524 32836 18528
rect 32772 18468 32776 18524
rect 32776 18468 32832 18524
rect 32832 18468 32836 18524
rect 32772 18464 32836 18468
rect 32852 18524 32916 18528
rect 32852 18468 32856 18524
rect 32856 18468 32912 18524
rect 32912 18468 32916 18524
rect 32852 18464 32916 18468
rect 37612 18524 37676 18528
rect 37612 18468 37616 18524
rect 37616 18468 37672 18524
rect 37672 18468 37676 18524
rect 37612 18464 37676 18468
rect 37692 18524 37756 18528
rect 37692 18468 37696 18524
rect 37696 18468 37752 18524
rect 37752 18468 37756 18524
rect 37692 18464 37756 18468
rect 37772 18524 37836 18528
rect 37772 18468 37776 18524
rect 37776 18468 37832 18524
rect 37832 18468 37836 18524
rect 37772 18464 37836 18468
rect 37852 18524 37916 18528
rect 37852 18468 37856 18524
rect 37856 18468 37912 18524
rect 37912 18468 37916 18524
rect 37852 18464 37916 18468
rect 1952 17980 2016 17984
rect 1952 17924 1956 17980
rect 1956 17924 2012 17980
rect 2012 17924 2016 17980
rect 1952 17920 2016 17924
rect 2032 17980 2096 17984
rect 2032 17924 2036 17980
rect 2036 17924 2092 17980
rect 2092 17924 2096 17980
rect 2032 17920 2096 17924
rect 2112 17980 2176 17984
rect 2112 17924 2116 17980
rect 2116 17924 2172 17980
rect 2172 17924 2176 17980
rect 2112 17920 2176 17924
rect 2192 17980 2256 17984
rect 2192 17924 2196 17980
rect 2196 17924 2252 17980
rect 2252 17924 2256 17980
rect 2192 17920 2256 17924
rect 6952 17980 7016 17984
rect 6952 17924 6956 17980
rect 6956 17924 7012 17980
rect 7012 17924 7016 17980
rect 6952 17920 7016 17924
rect 7032 17980 7096 17984
rect 7032 17924 7036 17980
rect 7036 17924 7092 17980
rect 7092 17924 7096 17980
rect 7032 17920 7096 17924
rect 7112 17980 7176 17984
rect 7112 17924 7116 17980
rect 7116 17924 7172 17980
rect 7172 17924 7176 17980
rect 7112 17920 7176 17924
rect 7192 17980 7256 17984
rect 7192 17924 7196 17980
rect 7196 17924 7252 17980
rect 7252 17924 7256 17980
rect 7192 17920 7256 17924
rect 11952 17980 12016 17984
rect 11952 17924 11956 17980
rect 11956 17924 12012 17980
rect 12012 17924 12016 17980
rect 11952 17920 12016 17924
rect 12032 17980 12096 17984
rect 12032 17924 12036 17980
rect 12036 17924 12092 17980
rect 12092 17924 12096 17980
rect 12032 17920 12096 17924
rect 12112 17980 12176 17984
rect 12112 17924 12116 17980
rect 12116 17924 12172 17980
rect 12172 17924 12176 17980
rect 12112 17920 12176 17924
rect 12192 17980 12256 17984
rect 12192 17924 12196 17980
rect 12196 17924 12252 17980
rect 12252 17924 12256 17980
rect 12192 17920 12256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 21952 17980 22016 17984
rect 21952 17924 21956 17980
rect 21956 17924 22012 17980
rect 22012 17924 22016 17980
rect 21952 17920 22016 17924
rect 22032 17980 22096 17984
rect 22032 17924 22036 17980
rect 22036 17924 22092 17980
rect 22092 17924 22096 17980
rect 22032 17920 22096 17924
rect 22112 17980 22176 17984
rect 22112 17924 22116 17980
rect 22116 17924 22172 17980
rect 22172 17924 22176 17980
rect 22112 17920 22176 17924
rect 22192 17980 22256 17984
rect 22192 17924 22196 17980
rect 22196 17924 22252 17980
rect 22252 17924 22256 17980
rect 22192 17920 22256 17924
rect 26952 17980 27016 17984
rect 26952 17924 26956 17980
rect 26956 17924 27012 17980
rect 27012 17924 27016 17980
rect 26952 17920 27016 17924
rect 27032 17980 27096 17984
rect 27032 17924 27036 17980
rect 27036 17924 27092 17980
rect 27092 17924 27096 17980
rect 27032 17920 27096 17924
rect 27112 17980 27176 17984
rect 27112 17924 27116 17980
rect 27116 17924 27172 17980
rect 27172 17924 27176 17980
rect 27112 17920 27176 17924
rect 27192 17980 27256 17984
rect 27192 17924 27196 17980
rect 27196 17924 27252 17980
rect 27252 17924 27256 17980
rect 27192 17920 27256 17924
rect 31952 17980 32016 17984
rect 31952 17924 31956 17980
rect 31956 17924 32012 17980
rect 32012 17924 32016 17980
rect 31952 17920 32016 17924
rect 32032 17980 32096 17984
rect 32032 17924 32036 17980
rect 32036 17924 32092 17980
rect 32092 17924 32096 17980
rect 32032 17920 32096 17924
rect 32112 17980 32176 17984
rect 32112 17924 32116 17980
rect 32116 17924 32172 17980
rect 32172 17924 32176 17980
rect 32112 17920 32176 17924
rect 32192 17980 32256 17984
rect 32192 17924 32196 17980
rect 32196 17924 32252 17980
rect 32252 17924 32256 17980
rect 32192 17920 32256 17924
rect 36952 17980 37016 17984
rect 36952 17924 36956 17980
rect 36956 17924 37012 17980
rect 37012 17924 37016 17980
rect 36952 17920 37016 17924
rect 37032 17980 37096 17984
rect 37032 17924 37036 17980
rect 37036 17924 37092 17980
rect 37092 17924 37096 17980
rect 37032 17920 37096 17924
rect 37112 17980 37176 17984
rect 37112 17924 37116 17980
rect 37116 17924 37172 17980
rect 37172 17924 37176 17980
rect 37112 17920 37176 17924
rect 37192 17980 37256 17984
rect 37192 17924 37196 17980
rect 37196 17924 37252 17980
rect 37252 17924 37256 17980
rect 37192 17920 37256 17924
rect 2612 17436 2676 17440
rect 2612 17380 2616 17436
rect 2616 17380 2672 17436
rect 2672 17380 2676 17436
rect 2612 17376 2676 17380
rect 2692 17436 2756 17440
rect 2692 17380 2696 17436
rect 2696 17380 2752 17436
rect 2752 17380 2756 17436
rect 2692 17376 2756 17380
rect 2772 17436 2836 17440
rect 2772 17380 2776 17436
rect 2776 17380 2832 17436
rect 2832 17380 2836 17436
rect 2772 17376 2836 17380
rect 2852 17436 2916 17440
rect 2852 17380 2856 17436
rect 2856 17380 2912 17436
rect 2912 17380 2916 17436
rect 2852 17376 2916 17380
rect 7612 17436 7676 17440
rect 7612 17380 7616 17436
rect 7616 17380 7672 17436
rect 7672 17380 7676 17436
rect 7612 17376 7676 17380
rect 7692 17436 7756 17440
rect 7692 17380 7696 17436
rect 7696 17380 7752 17436
rect 7752 17380 7756 17436
rect 7692 17376 7756 17380
rect 7772 17436 7836 17440
rect 7772 17380 7776 17436
rect 7776 17380 7832 17436
rect 7832 17380 7836 17436
rect 7772 17376 7836 17380
rect 7852 17436 7916 17440
rect 7852 17380 7856 17436
rect 7856 17380 7912 17436
rect 7912 17380 7916 17436
rect 7852 17376 7916 17380
rect 12612 17436 12676 17440
rect 12612 17380 12616 17436
rect 12616 17380 12672 17436
rect 12672 17380 12676 17436
rect 12612 17376 12676 17380
rect 12692 17436 12756 17440
rect 12692 17380 12696 17436
rect 12696 17380 12752 17436
rect 12752 17380 12756 17436
rect 12692 17376 12756 17380
rect 12772 17436 12836 17440
rect 12772 17380 12776 17436
rect 12776 17380 12832 17436
rect 12832 17380 12836 17436
rect 12772 17376 12836 17380
rect 12852 17436 12916 17440
rect 12852 17380 12856 17436
rect 12856 17380 12912 17436
rect 12912 17380 12916 17436
rect 12852 17376 12916 17380
rect 17612 17436 17676 17440
rect 17612 17380 17616 17436
rect 17616 17380 17672 17436
rect 17672 17380 17676 17436
rect 17612 17376 17676 17380
rect 17692 17436 17756 17440
rect 17692 17380 17696 17436
rect 17696 17380 17752 17436
rect 17752 17380 17756 17436
rect 17692 17376 17756 17380
rect 17772 17436 17836 17440
rect 17772 17380 17776 17436
rect 17776 17380 17832 17436
rect 17832 17380 17836 17436
rect 17772 17376 17836 17380
rect 17852 17436 17916 17440
rect 17852 17380 17856 17436
rect 17856 17380 17912 17436
rect 17912 17380 17916 17436
rect 17852 17376 17916 17380
rect 22612 17436 22676 17440
rect 22612 17380 22616 17436
rect 22616 17380 22672 17436
rect 22672 17380 22676 17436
rect 22612 17376 22676 17380
rect 22692 17436 22756 17440
rect 22692 17380 22696 17436
rect 22696 17380 22752 17436
rect 22752 17380 22756 17436
rect 22692 17376 22756 17380
rect 22772 17436 22836 17440
rect 22772 17380 22776 17436
rect 22776 17380 22832 17436
rect 22832 17380 22836 17436
rect 22772 17376 22836 17380
rect 22852 17436 22916 17440
rect 22852 17380 22856 17436
rect 22856 17380 22912 17436
rect 22912 17380 22916 17436
rect 22852 17376 22916 17380
rect 27612 17436 27676 17440
rect 27612 17380 27616 17436
rect 27616 17380 27672 17436
rect 27672 17380 27676 17436
rect 27612 17376 27676 17380
rect 27692 17436 27756 17440
rect 27692 17380 27696 17436
rect 27696 17380 27752 17436
rect 27752 17380 27756 17436
rect 27692 17376 27756 17380
rect 27772 17436 27836 17440
rect 27772 17380 27776 17436
rect 27776 17380 27832 17436
rect 27832 17380 27836 17436
rect 27772 17376 27836 17380
rect 27852 17436 27916 17440
rect 27852 17380 27856 17436
rect 27856 17380 27912 17436
rect 27912 17380 27916 17436
rect 27852 17376 27916 17380
rect 32612 17436 32676 17440
rect 32612 17380 32616 17436
rect 32616 17380 32672 17436
rect 32672 17380 32676 17436
rect 32612 17376 32676 17380
rect 32692 17436 32756 17440
rect 32692 17380 32696 17436
rect 32696 17380 32752 17436
rect 32752 17380 32756 17436
rect 32692 17376 32756 17380
rect 32772 17436 32836 17440
rect 32772 17380 32776 17436
rect 32776 17380 32832 17436
rect 32832 17380 32836 17436
rect 32772 17376 32836 17380
rect 32852 17436 32916 17440
rect 32852 17380 32856 17436
rect 32856 17380 32912 17436
rect 32912 17380 32916 17436
rect 32852 17376 32916 17380
rect 37612 17436 37676 17440
rect 37612 17380 37616 17436
rect 37616 17380 37672 17436
rect 37672 17380 37676 17436
rect 37612 17376 37676 17380
rect 37692 17436 37756 17440
rect 37692 17380 37696 17436
rect 37696 17380 37752 17436
rect 37752 17380 37756 17436
rect 37692 17376 37756 17380
rect 37772 17436 37836 17440
rect 37772 17380 37776 17436
rect 37776 17380 37832 17436
rect 37832 17380 37836 17436
rect 37772 17376 37836 17380
rect 37852 17436 37916 17440
rect 37852 17380 37856 17436
rect 37856 17380 37912 17436
rect 37912 17380 37916 17436
rect 37852 17376 37916 17380
rect 1952 16892 2016 16896
rect 1952 16836 1956 16892
rect 1956 16836 2012 16892
rect 2012 16836 2016 16892
rect 1952 16832 2016 16836
rect 2032 16892 2096 16896
rect 2032 16836 2036 16892
rect 2036 16836 2092 16892
rect 2092 16836 2096 16892
rect 2032 16832 2096 16836
rect 2112 16892 2176 16896
rect 2112 16836 2116 16892
rect 2116 16836 2172 16892
rect 2172 16836 2176 16892
rect 2112 16832 2176 16836
rect 2192 16892 2256 16896
rect 2192 16836 2196 16892
rect 2196 16836 2252 16892
rect 2252 16836 2256 16892
rect 2192 16832 2256 16836
rect 6952 16892 7016 16896
rect 6952 16836 6956 16892
rect 6956 16836 7012 16892
rect 7012 16836 7016 16892
rect 6952 16832 7016 16836
rect 7032 16892 7096 16896
rect 7032 16836 7036 16892
rect 7036 16836 7092 16892
rect 7092 16836 7096 16892
rect 7032 16832 7096 16836
rect 7112 16892 7176 16896
rect 7112 16836 7116 16892
rect 7116 16836 7172 16892
rect 7172 16836 7176 16892
rect 7112 16832 7176 16836
rect 7192 16892 7256 16896
rect 7192 16836 7196 16892
rect 7196 16836 7252 16892
rect 7252 16836 7256 16892
rect 7192 16832 7256 16836
rect 11952 16892 12016 16896
rect 11952 16836 11956 16892
rect 11956 16836 12012 16892
rect 12012 16836 12016 16892
rect 11952 16832 12016 16836
rect 12032 16892 12096 16896
rect 12032 16836 12036 16892
rect 12036 16836 12092 16892
rect 12092 16836 12096 16892
rect 12032 16832 12096 16836
rect 12112 16892 12176 16896
rect 12112 16836 12116 16892
rect 12116 16836 12172 16892
rect 12172 16836 12176 16892
rect 12112 16832 12176 16836
rect 12192 16892 12256 16896
rect 12192 16836 12196 16892
rect 12196 16836 12252 16892
rect 12252 16836 12256 16892
rect 12192 16832 12256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 21952 16892 22016 16896
rect 21952 16836 21956 16892
rect 21956 16836 22012 16892
rect 22012 16836 22016 16892
rect 21952 16832 22016 16836
rect 22032 16892 22096 16896
rect 22032 16836 22036 16892
rect 22036 16836 22092 16892
rect 22092 16836 22096 16892
rect 22032 16832 22096 16836
rect 22112 16892 22176 16896
rect 22112 16836 22116 16892
rect 22116 16836 22172 16892
rect 22172 16836 22176 16892
rect 22112 16832 22176 16836
rect 22192 16892 22256 16896
rect 22192 16836 22196 16892
rect 22196 16836 22252 16892
rect 22252 16836 22256 16892
rect 22192 16832 22256 16836
rect 26952 16892 27016 16896
rect 26952 16836 26956 16892
rect 26956 16836 27012 16892
rect 27012 16836 27016 16892
rect 26952 16832 27016 16836
rect 27032 16892 27096 16896
rect 27032 16836 27036 16892
rect 27036 16836 27092 16892
rect 27092 16836 27096 16892
rect 27032 16832 27096 16836
rect 27112 16892 27176 16896
rect 27112 16836 27116 16892
rect 27116 16836 27172 16892
rect 27172 16836 27176 16892
rect 27112 16832 27176 16836
rect 27192 16892 27256 16896
rect 27192 16836 27196 16892
rect 27196 16836 27252 16892
rect 27252 16836 27256 16892
rect 27192 16832 27256 16836
rect 31952 16892 32016 16896
rect 31952 16836 31956 16892
rect 31956 16836 32012 16892
rect 32012 16836 32016 16892
rect 31952 16832 32016 16836
rect 32032 16892 32096 16896
rect 32032 16836 32036 16892
rect 32036 16836 32092 16892
rect 32092 16836 32096 16892
rect 32032 16832 32096 16836
rect 32112 16892 32176 16896
rect 32112 16836 32116 16892
rect 32116 16836 32172 16892
rect 32172 16836 32176 16892
rect 32112 16832 32176 16836
rect 32192 16892 32256 16896
rect 32192 16836 32196 16892
rect 32196 16836 32252 16892
rect 32252 16836 32256 16892
rect 32192 16832 32256 16836
rect 36952 16892 37016 16896
rect 36952 16836 36956 16892
rect 36956 16836 37012 16892
rect 37012 16836 37016 16892
rect 36952 16832 37016 16836
rect 37032 16892 37096 16896
rect 37032 16836 37036 16892
rect 37036 16836 37092 16892
rect 37092 16836 37096 16892
rect 37032 16832 37096 16836
rect 37112 16892 37176 16896
rect 37112 16836 37116 16892
rect 37116 16836 37172 16892
rect 37172 16836 37176 16892
rect 37112 16832 37176 16836
rect 37192 16892 37256 16896
rect 37192 16836 37196 16892
rect 37196 16836 37252 16892
rect 37252 16836 37256 16892
rect 37192 16832 37256 16836
rect 2612 16348 2676 16352
rect 2612 16292 2616 16348
rect 2616 16292 2672 16348
rect 2672 16292 2676 16348
rect 2612 16288 2676 16292
rect 2692 16348 2756 16352
rect 2692 16292 2696 16348
rect 2696 16292 2752 16348
rect 2752 16292 2756 16348
rect 2692 16288 2756 16292
rect 2772 16348 2836 16352
rect 2772 16292 2776 16348
rect 2776 16292 2832 16348
rect 2832 16292 2836 16348
rect 2772 16288 2836 16292
rect 2852 16348 2916 16352
rect 2852 16292 2856 16348
rect 2856 16292 2912 16348
rect 2912 16292 2916 16348
rect 2852 16288 2916 16292
rect 7612 16348 7676 16352
rect 7612 16292 7616 16348
rect 7616 16292 7672 16348
rect 7672 16292 7676 16348
rect 7612 16288 7676 16292
rect 7692 16348 7756 16352
rect 7692 16292 7696 16348
rect 7696 16292 7752 16348
rect 7752 16292 7756 16348
rect 7692 16288 7756 16292
rect 7772 16348 7836 16352
rect 7772 16292 7776 16348
rect 7776 16292 7832 16348
rect 7832 16292 7836 16348
rect 7772 16288 7836 16292
rect 7852 16348 7916 16352
rect 7852 16292 7856 16348
rect 7856 16292 7912 16348
rect 7912 16292 7916 16348
rect 7852 16288 7916 16292
rect 12612 16348 12676 16352
rect 12612 16292 12616 16348
rect 12616 16292 12672 16348
rect 12672 16292 12676 16348
rect 12612 16288 12676 16292
rect 12692 16348 12756 16352
rect 12692 16292 12696 16348
rect 12696 16292 12752 16348
rect 12752 16292 12756 16348
rect 12692 16288 12756 16292
rect 12772 16348 12836 16352
rect 12772 16292 12776 16348
rect 12776 16292 12832 16348
rect 12832 16292 12836 16348
rect 12772 16288 12836 16292
rect 12852 16348 12916 16352
rect 12852 16292 12856 16348
rect 12856 16292 12912 16348
rect 12912 16292 12916 16348
rect 12852 16288 12916 16292
rect 17612 16348 17676 16352
rect 17612 16292 17616 16348
rect 17616 16292 17672 16348
rect 17672 16292 17676 16348
rect 17612 16288 17676 16292
rect 17692 16348 17756 16352
rect 17692 16292 17696 16348
rect 17696 16292 17752 16348
rect 17752 16292 17756 16348
rect 17692 16288 17756 16292
rect 17772 16348 17836 16352
rect 17772 16292 17776 16348
rect 17776 16292 17832 16348
rect 17832 16292 17836 16348
rect 17772 16288 17836 16292
rect 17852 16348 17916 16352
rect 17852 16292 17856 16348
rect 17856 16292 17912 16348
rect 17912 16292 17916 16348
rect 17852 16288 17916 16292
rect 22612 16348 22676 16352
rect 22612 16292 22616 16348
rect 22616 16292 22672 16348
rect 22672 16292 22676 16348
rect 22612 16288 22676 16292
rect 22692 16348 22756 16352
rect 22692 16292 22696 16348
rect 22696 16292 22752 16348
rect 22752 16292 22756 16348
rect 22692 16288 22756 16292
rect 22772 16348 22836 16352
rect 22772 16292 22776 16348
rect 22776 16292 22832 16348
rect 22832 16292 22836 16348
rect 22772 16288 22836 16292
rect 22852 16348 22916 16352
rect 22852 16292 22856 16348
rect 22856 16292 22912 16348
rect 22912 16292 22916 16348
rect 22852 16288 22916 16292
rect 27612 16348 27676 16352
rect 27612 16292 27616 16348
rect 27616 16292 27672 16348
rect 27672 16292 27676 16348
rect 27612 16288 27676 16292
rect 27692 16348 27756 16352
rect 27692 16292 27696 16348
rect 27696 16292 27752 16348
rect 27752 16292 27756 16348
rect 27692 16288 27756 16292
rect 27772 16348 27836 16352
rect 27772 16292 27776 16348
rect 27776 16292 27832 16348
rect 27832 16292 27836 16348
rect 27772 16288 27836 16292
rect 27852 16348 27916 16352
rect 27852 16292 27856 16348
rect 27856 16292 27912 16348
rect 27912 16292 27916 16348
rect 27852 16288 27916 16292
rect 32612 16348 32676 16352
rect 32612 16292 32616 16348
rect 32616 16292 32672 16348
rect 32672 16292 32676 16348
rect 32612 16288 32676 16292
rect 32692 16348 32756 16352
rect 32692 16292 32696 16348
rect 32696 16292 32752 16348
rect 32752 16292 32756 16348
rect 32692 16288 32756 16292
rect 32772 16348 32836 16352
rect 32772 16292 32776 16348
rect 32776 16292 32832 16348
rect 32832 16292 32836 16348
rect 32772 16288 32836 16292
rect 32852 16348 32916 16352
rect 32852 16292 32856 16348
rect 32856 16292 32912 16348
rect 32912 16292 32916 16348
rect 32852 16288 32916 16292
rect 37612 16348 37676 16352
rect 37612 16292 37616 16348
rect 37616 16292 37672 16348
rect 37672 16292 37676 16348
rect 37612 16288 37676 16292
rect 37692 16348 37756 16352
rect 37692 16292 37696 16348
rect 37696 16292 37752 16348
rect 37752 16292 37756 16348
rect 37692 16288 37756 16292
rect 37772 16348 37836 16352
rect 37772 16292 37776 16348
rect 37776 16292 37832 16348
rect 37832 16292 37836 16348
rect 37772 16288 37836 16292
rect 37852 16348 37916 16352
rect 37852 16292 37856 16348
rect 37856 16292 37912 16348
rect 37912 16292 37916 16348
rect 37852 16288 37916 16292
rect 1952 15804 2016 15808
rect 1952 15748 1956 15804
rect 1956 15748 2012 15804
rect 2012 15748 2016 15804
rect 1952 15744 2016 15748
rect 2032 15804 2096 15808
rect 2032 15748 2036 15804
rect 2036 15748 2092 15804
rect 2092 15748 2096 15804
rect 2032 15744 2096 15748
rect 2112 15804 2176 15808
rect 2112 15748 2116 15804
rect 2116 15748 2172 15804
rect 2172 15748 2176 15804
rect 2112 15744 2176 15748
rect 2192 15804 2256 15808
rect 2192 15748 2196 15804
rect 2196 15748 2252 15804
rect 2252 15748 2256 15804
rect 2192 15744 2256 15748
rect 6952 15804 7016 15808
rect 6952 15748 6956 15804
rect 6956 15748 7012 15804
rect 7012 15748 7016 15804
rect 6952 15744 7016 15748
rect 7032 15804 7096 15808
rect 7032 15748 7036 15804
rect 7036 15748 7092 15804
rect 7092 15748 7096 15804
rect 7032 15744 7096 15748
rect 7112 15804 7176 15808
rect 7112 15748 7116 15804
rect 7116 15748 7172 15804
rect 7172 15748 7176 15804
rect 7112 15744 7176 15748
rect 7192 15804 7256 15808
rect 7192 15748 7196 15804
rect 7196 15748 7252 15804
rect 7252 15748 7256 15804
rect 7192 15744 7256 15748
rect 11952 15804 12016 15808
rect 11952 15748 11956 15804
rect 11956 15748 12012 15804
rect 12012 15748 12016 15804
rect 11952 15744 12016 15748
rect 12032 15804 12096 15808
rect 12032 15748 12036 15804
rect 12036 15748 12092 15804
rect 12092 15748 12096 15804
rect 12032 15744 12096 15748
rect 12112 15804 12176 15808
rect 12112 15748 12116 15804
rect 12116 15748 12172 15804
rect 12172 15748 12176 15804
rect 12112 15744 12176 15748
rect 12192 15804 12256 15808
rect 12192 15748 12196 15804
rect 12196 15748 12252 15804
rect 12252 15748 12256 15804
rect 12192 15744 12256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 21952 15804 22016 15808
rect 21952 15748 21956 15804
rect 21956 15748 22012 15804
rect 22012 15748 22016 15804
rect 21952 15744 22016 15748
rect 22032 15804 22096 15808
rect 22032 15748 22036 15804
rect 22036 15748 22092 15804
rect 22092 15748 22096 15804
rect 22032 15744 22096 15748
rect 22112 15804 22176 15808
rect 22112 15748 22116 15804
rect 22116 15748 22172 15804
rect 22172 15748 22176 15804
rect 22112 15744 22176 15748
rect 22192 15804 22256 15808
rect 22192 15748 22196 15804
rect 22196 15748 22252 15804
rect 22252 15748 22256 15804
rect 22192 15744 22256 15748
rect 26952 15804 27016 15808
rect 26952 15748 26956 15804
rect 26956 15748 27012 15804
rect 27012 15748 27016 15804
rect 26952 15744 27016 15748
rect 27032 15804 27096 15808
rect 27032 15748 27036 15804
rect 27036 15748 27092 15804
rect 27092 15748 27096 15804
rect 27032 15744 27096 15748
rect 27112 15804 27176 15808
rect 27112 15748 27116 15804
rect 27116 15748 27172 15804
rect 27172 15748 27176 15804
rect 27112 15744 27176 15748
rect 27192 15804 27256 15808
rect 27192 15748 27196 15804
rect 27196 15748 27252 15804
rect 27252 15748 27256 15804
rect 27192 15744 27256 15748
rect 31952 15804 32016 15808
rect 31952 15748 31956 15804
rect 31956 15748 32012 15804
rect 32012 15748 32016 15804
rect 31952 15744 32016 15748
rect 32032 15804 32096 15808
rect 32032 15748 32036 15804
rect 32036 15748 32092 15804
rect 32092 15748 32096 15804
rect 32032 15744 32096 15748
rect 32112 15804 32176 15808
rect 32112 15748 32116 15804
rect 32116 15748 32172 15804
rect 32172 15748 32176 15804
rect 32112 15744 32176 15748
rect 32192 15804 32256 15808
rect 32192 15748 32196 15804
rect 32196 15748 32252 15804
rect 32252 15748 32256 15804
rect 32192 15744 32256 15748
rect 36952 15804 37016 15808
rect 36952 15748 36956 15804
rect 36956 15748 37012 15804
rect 37012 15748 37016 15804
rect 36952 15744 37016 15748
rect 37032 15804 37096 15808
rect 37032 15748 37036 15804
rect 37036 15748 37092 15804
rect 37092 15748 37096 15804
rect 37032 15744 37096 15748
rect 37112 15804 37176 15808
rect 37112 15748 37116 15804
rect 37116 15748 37172 15804
rect 37172 15748 37176 15804
rect 37112 15744 37176 15748
rect 37192 15804 37256 15808
rect 37192 15748 37196 15804
rect 37196 15748 37252 15804
rect 37252 15748 37256 15804
rect 37192 15744 37256 15748
rect 2612 15260 2676 15264
rect 2612 15204 2616 15260
rect 2616 15204 2672 15260
rect 2672 15204 2676 15260
rect 2612 15200 2676 15204
rect 2692 15260 2756 15264
rect 2692 15204 2696 15260
rect 2696 15204 2752 15260
rect 2752 15204 2756 15260
rect 2692 15200 2756 15204
rect 2772 15260 2836 15264
rect 2772 15204 2776 15260
rect 2776 15204 2832 15260
rect 2832 15204 2836 15260
rect 2772 15200 2836 15204
rect 2852 15260 2916 15264
rect 2852 15204 2856 15260
rect 2856 15204 2912 15260
rect 2912 15204 2916 15260
rect 2852 15200 2916 15204
rect 7612 15260 7676 15264
rect 7612 15204 7616 15260
rect 7616 15204 7672 15260
rect 7672 15204 7676 15260
rect 7612 15200 7676 15204
rect 7692 15260 7756 15264
rect 7692 15204 7696 15260
rect 7696 15204 7752 15260
rect 7752 15204 7756 15260
rect 7692 15200 7756 15204
rect 7772 15260 7836 15264
rect 7772 15204 7776 15260
rect 7776 15204 7832 15260
rect 7832 15204 7836 15260
rect 7772 15200 7836 15204
rect 7852 15260 7916 15264
rect 7852 15204 7856 15260
rect 7856 15204 7912 15260
rect 7912 15204 7916 15260
rect 7852 15200 7916 15204
rect 12612 15260 12676 15264
rect 12612 15204 12616 15260
rect 12616 15204 12672 15260
rect 12672 15204 12676 15260
rect 12612 15200 12676 15204
rect 12692 15260 12756 15264
rect 12692 15204 12696 15260
rect 12696 15204 12752 15260
rect 12752 15204 12756 15260
rect 12692 15200 12756 15204
rect 12772 15260 12836 15264
rect 12772 15204 12776 15260
rect 12776 15204 12832 15260
rect 12832 15204 12836 15260
rect 12772 15200 12836 15204
rect 12852 15260 12916 15264
rect 12852 15204 12856 15260
rect 12856 15204 12912 15260
rect 12912 15204 12916 15260
rect 12852 15200 12916 15204
rect 17612 15260 17676 15264
rect 17612 15204 17616 15260
rect 17616 15204 17672 15260
rect 17672 15204 17676 15260
rect 17612 15200 17676 15204
rect 17692 15260 17756 15264
rect 17692 15204 17696 15260
rect 17696 15204 17752 15260
rect 17752 15204 17756 15260
rect 17692 15200 17756 15204
rect 17772 15260 17836 15264
rect 17772 15204 17776 15260
rect 17776 15204 17832 15260
rect 17832 15204 17836 15260
rect 17772 15200 17836 15204
rect 17852 15260 17916 15264
rect 17852 15204 17856 15260
rect 17856 15204 17912 15260
rect 17912 15204 17916 15260
rect 17852 15200 17916 15204
rect 22612 15260 22676 15264
rect 22612 15204 22616 15260
rect 22616 15204 22672 15260
rect 22672 15204 22676 15260
rect 22612 15200 22676 15204
rect 22692 15260 22756 15264
rect 22692 15204 22696 15260
rect 22696 15204 22752 15260
rect 22752 15204 22756 15260
rect 22692 15200 22756 15204
rect 22772 15260 22836 15264
rect 22772 15204 22776 15260
rect 22776 15204 22832 15260
rect 22832 15204 22836 15260
rect 22772 15200 22836 15204
rect 22852 15260 22916 15264
rect 22852 15204 22856 15260
rect 22856 15204 22912 15260
rect 22912 15204 22916 15260
rect 22852 15200 22916 15204
rect 27612 15260 27676 15264
rect 27612 15204 27616 15260
rect 27616 15204 27672 15260
rect 27672 15204 27676 15260
rect 27612 15200 27676 15204
rect 27692 15260 27756 15264
rect 27692 15204 27696 15260
rect 27696 15204 27752 15260
rect 27752 15204 27756 15260
rect 27692 15200 27756 15204
rect 27772 15260 27836 15264
rect 27772 15204 27776 15260
rect 27776 15204 27832 15260
rect 27832 15204 27836 15260
rect 27772 15200 27836 15204
rect 27852 15260 27916 15264
rect 27852 15204 27856 15260
rect 27856 15204 27912 15260
rect 27912 15204 27916 15260
rect 27852 15200 27916 15204
rect 32612 15260 32676 15264
rect 32612 15204 32616 15260
rect 32616 15204 32672 15260
rect 32672 15204 32676 15260
rect 32612 15200 32676 15204
rect 32692 15260 32756 15264
rect 32692 15204 32696 15260
rect 32696 15204 32752 15260
rect 32752 15204 32756 15260
rect 32692 15200 32756 15204
rect 32772 15260 32836 15264
rect 32772 15204 32776 15260
rect 32776 15204 32832 15260
rect 32832 15204 32836 15260
rect 32772 15200 32836 15204
rect 32852 15260 32916 15264
rect 32852 15204 32856 15260
rect 32856 15204 32912 15260
rect 32912 15204 32916 15260
rect 32852 15200 32916 15204
rect 37612 15260 37676 15264
rect 37612 15204 37616 15260
rect 37616 15204 37672 15260
rect 37672 15204 37676 15260
rect 37612 15200 37676 15204
rect 37692 15260 37756 15264
rect 37692 15204 37696 15260
rect 37696 15204 37752 15260
rect 37752 15204 37756 15260
rect 37692 15200 37756 15204
rect 37772 15260 37836 15264
rect 37772 15204 37776 15260
rect 37776 15204 37832 15260
rect 37832 15204 37836 15260
rect 37772 15200 37836 15204
rect 37852 15260 37916 15264
rect 37852 15204 37856 15260
rect 37856 15204 37912 15260
rect 37912 15204 37916 15260
rect 37852 15200 37916 15204
rect 1952 14716 2016 14720
rect 1952 14660 1956 14716
rect 1956 14660 2012 14716
rect 2012 14660 2016 14716
rect 1952 14656 2016 14660
rect 2032 14716 2096 14720
rect 2032 14660 2036 14716
rect 2036 14660 2092 14716
rect 2092 14660 2096 14716
rect 2032 14656 2096 14660
rect 2112 14716 2176 14720
rect 2112 14660 2116 14716
rect 2116 14660 2172 14716
rect 2172 14660 2176 14716
rect 2112 14656 2176 14660
rect 2192 14716 2256 14720
rect 2192 14660 2196 14716
rect 2196 14660 2252 14716
rect 2252 14660 2256 14716
rect 2192 14656 2256 14660
rect 6952 14716 7016 14720
rect 6952 14660 6956 14716
rect 6956 14660 7012 14716
rect 7012 14660 7016 14716
rect 6952 14656 7016 14660
rect 7032 14716 7096 14720
rect 7032 14660 7036 14716
rect 7036 14660 7092 14716
rect 7092 14660 7096 14716
rect 7032 14656 7096 14660
rect 7112 14716 7176 14720
rect 7112 14660 7116 14716
rect 7116 14660 7172 14716
rect 7172 14660 7176 14716
rect 7112 14656 7176 14660
rect 7192 14716 7256 14720
rect 7192 14660 7196 14716
rect 7196 14660 7252 14716
rect 7252 14660 7256 14716
rect 7192 14656 7256 14660
rect 11952 14716 12016 14720
rect 11952 14660 11956 14716
rect 11956 14660 12012 14716
rect 12012 14660 12016 14716
rect 11952 14656 12016 14660
rect 12032 14716 12096 14720
rect 12032 14660 12036 14716
rect 12036 14660 12092 14716
rect 12092 14660 12096 14716
rect 12032 14656 12096 14660
rect 12112 14716 12176 14720
rect 12112 14660 12116 14716
rect 12116 14660 12172 14716
rect 12172 14660 12176 14716
rect 12112 14656 12176 14660
rect 12192 14716 12256 14720
rect 12192 14660 12196 14716
rect 12196 14660 12252 14716
rect 12252 14660 12256 14716
rect 12192 14656 12256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 21952 14716 22016 14720
rect 21952 14660 21956 14716
rect 21956 14660 22012 14716
rect 22012 14660 22016 14716
rect 21952 14656 22016 14660
rect 22032 14716 22096 14720
rect 22032 14660 22036 14716
rect 22036 14660 22092 14716
rect 22092 14660 22096 14716
rect 22032 14656 22096 14660
rect 22112 14716 22176 14720
rect 22112 14660 22116 14716
rect 22116 14660 22172 14716
rect 22172 14660 22176 14716
rect 22112 14656 22176 14660
rect 22192 14716 22256 14720
rect 22192 14660 22196 14716
rect 22196 14660 22252 14716
rect 22252 14660 22256 14716
rect 22192 14656 22256 14660
rect 26952 14716 27016 14720
rect 26952 14660 26956 14716
rect 26956 14660 27012 14716
rect 27012 14660 27016 14716
rect 26952 14656 27016 14660
rect 27032 14716 27096 14720
rect 27032 14660 27036 14716
rect 27036 14660 27092 14716
rect 27092 14660 27096 14716
rect 27032 14656 27096 14660
rect 27112 14716 27176 14720
rect 27112 14660 27116 14716
rect 27116 14660 27172 14716
rect 27172 14660 27176 14716
rect 27112 14656 27176 14660
rect 27192 14716 27256 14720
rect 27192 14660 27196 14716
rect 27196 14660 27252 14716
rect 27252 14660 27256 14716
rect 27192 14656 27256 14660
rect 31952 14716 32016 14720
rect 31952 14660 31956 14716
rect 31956 14660 32012 14716
rect 32012 14660 32016 14716
rect 31952 14656 32016 14660
rect 32032 14716 32096 14720
rect 32032 14660 32036 14716
rect 32036 14660 32092 14716
rect 32092 14660 32096 14716
rect 32032 14656 32096 14660
rect 32112 14716 32176 14720
rect 32112 14660 32116 14716
rect 32116 14660 32172 14716
rect 32172 14660 32176 14716
rect 32112 14656 32176 14660
rect 32192 14716 32256 14720
rect 32192 14660 32196 14716
rect 32196 14660 32252 14716
rect 32252 14660 32256 14716
rect 32192 14656 32256 14660
rect 36952 14716 37016 14720
rect 36952 14660 36956 14716
rect 36956 14660 37012 14716
rect 37012 14660 37016 14716
rect 36952 14656 37016 14660
rect 37032 14716 37096 14720
rect 37032 14660 37036 14716
rect 37036 14660 37092 14716
rect 37092 14660 37096 14716
rect 37032 14656 37096 14660
rect 37112 14716 37176 14720
rect 37112 14660 37116 14716
rect 37116 14660 37172 14716
rect 37172 14660 37176 14716
rect 37112 14656 37176 14660
rect 37192 14716 37256 14720
rect 37192 14660 37196 14716
rect 37196 14660 37252 14716
rect 37252 14660 37256 14716
rect 37192 14656 37256 14660
rect 2612 14172 2676 14176
rect 2612 14116 2616 14172
rect 2616 14116 2672 14172
rect 2672 14116 2676 14172
rect 2612 14112 2676 14116
rect 2692 14172 2756 14176
rect 2692 14116 2696 14172
rect 2696 14116 2752 14172
rect 2752 14116 2756 14172
rect 2692 14112 2756 14116
rect 2772 14172 2836 14176
rect 2772 14116 2776 14172
rect 2776 14116 2832 14172
rect 2832 14116 2836 14172
rect 2772 14112 2836 14116
rect 2852 14172 2916 14176
rect 2852 14116 2856 14172
rect 2856 14116 2912 14172
rect 2912 14116 2916 14172
rect 2852 14112 2916 14116
rect 7612 14172 7676 14176
rect 7612 14116 7616 14172
rect 7616 14116 7672 14172
rect 7672 14116 7676 14172
rect 7612 14112 7676 14116
rect 7692 14172 7756 14176
rect 7692 14116 7696 14172
rect 7696 14116 7752 14172
rect 7752 14116 7756 14172
rect 7692 14112 7756 14116
rect 7772 14172 7836 14176
rect 7772 14116 7776 14172
rect 7776 14116 7832 14172
rect 7832 14116 7836 14172
rect 7772 14112 7836 14116
rect 7852 14172 7916 14176
rect 7852 14116 7856 14172
rect 7856 14116 7912 14172
rect 7912 14116 7916 14172
rect 7852 14112 7916 14116
rect 12612 14172 12676 14176
rect 12612 14116 12616 14172
rect 12616 14116 12672 14172
rect 12672 14116 12676 14172
rect 12612 14112 12676 14116
rect 12692 14172 12756 14176
rect 12692 14116 12696 14172
rect 12696 14116 12752 14172
rect 12752 14116 12756 14172
rect 12692 14112 12756 14116
rect 12772 14172 12836 14176
rect 12772 14116 12776 14172
rect 12776 14116 12832 14172
rect 12832 14116 12836 14172
rect 12772 14112 12836 14116
rect 12852 14172 12916 14176
rect 12852 14116 12856 14172
rect 12856 14116 12912 14172
rect 12912 14116 12916 14172
rect 12852 14112 12916 14116
rect 17612 14172 17676 14176
rect 17612 14116 17616 14172
rect 17616 14116 17672 14172
rect 17672 14116 17676 14172
rect 17612 14112 17676 14116
rect 17692 14172 17756 14176
rect 17692 14116 17696 14172
rect 17696 14116 17752 14172
rect 17752 14116 17756 14172
rect 17692 14112 17756 14116
rect 17772 14172 17836 14176
rect 17772 14116 17776 14172
rect 17776 14116 17832 14172
rect 17832 14116 17836 14172
rect 17772 14112 17836 14116
rect 17852 14172 17916 14176
rect 17852 14116 17856 14172
rect 17856 14116 17912 14172
rect 17912 14116 17916 14172
rect 17852 14112 17916 14116
rect 22612 14172 22676 14176
rect 22612 14116 22616 14172
rect 22616 14116 22672 14172
rect 22672 14116 22676 14172
rect 22612 14112 22676 14116
rect 22692 14172 22756 14176
rect 22692 14116 22696 14172
rect 22696 14116 22752 14172
rect 22752 14116 22756 14172
rect 22692 14112 22756 14116
rect 22772 14172 22836 14176
rect 22772 14116 22776 14172
rect 22776 14116 22832 14172
rect 22832 14116 22836 14172
rect 22772 14112 22836 14116
rect 22852 14172 22916 14176
rect 22852 14116 22856 14172
rect 22856 14116 22912 14172
rect 22912 14116 22916 14172
rect 22852 14112 22916 14116
rect 27612 14172 27676 14176
rect 27612 14116 27616 14172
rect 27616 14116 27672 14172
rect 27672 14116 27676 14172
rect 27612 14112 27676 14116
rect 27692 14172 27756 14176
rect 27692 14116 27696 14172
rect 27696 14116 27752 14172
rect 27752 14116 27756 14172
rect 27692 14112 27756 14116
rect 27772 14172 27836 14176
rect 27772 14116 27776 14172
rect 27776 14116 27832 14172
rect 27832 14116 27836 14172
rect 27772 14112 27836 14116
rect 27852 14172 27916 14176
rect 27852 14116 27856 14172
rect 27856 14116 27912 14172
rect 27912 14116 27916 14172
rect 27852 14112 27916 14116
rect 32612 14172 32676 14176
rect 32612 14116 32616 14172
rect 32616 14116 32672 14172
rect 32672 14116 32676 14172
rect 32612 14112 32676 14116
rect 32692 14172 32756 14176
rect 32692 14116 32696 14172
rect 32696 14116 32752 14172
rect 32752 14116 32756 14172
rect 32692 14112 32756 14116
rect 32772 14172 32836 14176
rect 32772 14116 32776 14172
rect 32776 14116 32832 14172
rect 32832 14116 32836 14172
rect 32772 14112 32836 14116
rect 32852 14172 32916 14176
rect 32852 14116 32856 14172
rect 32856 14116 32912 14172
rect 32912 14116 32916 14172
rect 32852 14112 32916 14116
rect 37612 14172 37676 14176
rect 37612 14116 37616 14172
rect 37616 14116 37672 14172
rect 37672 14116 37676 14172
rect 37612 14112 37676 14116
rect 37692 14172 37756 14176
rect 37692 14116 37696 14172
rect 37696 14116 37752 14172
rect 37752 14116 37756 14172
rect 37692 14112 37756 14116
rect 37772 14172 37836 14176
rect 37772 14116 37776 14172
rect 37776 14116 37832 14172
rect 37832 14116 37836 14172
rect 37772 14112 37836 14116
rect 37852 14172 37916 14176
rect 37852 14116 37856 14172
rect 37856 14116 37912 14172
rect 37912 14116 37916 14172
rect 37852 14112 37916 14116
rect 1952 13628 2016 13632
rect 1952 13572 1956 13628
rect 1956 13572 2012 13628
rect 2012 13572 2016 13628
rect 1952 13568 2016 13572
rect 2032 13628 2096 13632
rect 2032 13572 2036 13628
rect 2036 13572 2092 13628
rect 2092 13572 2096 13628
rect 2032 13568 2096 13572
rect 2112 13628 2176 13632
rect 2112 13572 2116 13628
rect 2116 13572 2172 13628
rect 2172 13572 2176 13628
rect 2112 13568 2176 13572
rect 2192 13628 2256 13632
rect 2192 13572 2196 13628
rect 2196 13572 2252 13628
rect 2252 13572 2256 13628
rect 2192 13568 2256 13572
rect 6952 13628 7016 13632
rect 6952 13572 6956 13628
rect 6956 13572 7012 13628
rect 7012 13572 7016 13628
rect 6952 13568 7016 13572
rect 7032 13628 7096 13632
rect 7032 13572 7036 13628
rect 7036 13572 7092 13628
rect 7092 13572 7096 13628
rect 7032 13568 7096 13572
rect 7112 13628 7176 13632
rect 7112 13572 7116 13628
rect 7116 13572 7172 13628
rect 7172 13572 7176 13628
rect 7112 13568 7176 13572
rect 7192 13628 7256 13632
rect 7192 13572 7196 13628
rect 7196 13572 7252 13628
rect 7252 13572 7256 13628
rect 7192 13568 7256 13572
rect 11952 13628 12016 13632
rect 11952 13572 11956 13628
rect 11956 13572 12012 13628
rect 12012 13572 12016 13628
rect 11952 13568 12016 13572
rect 12032 13628 12096 13632
rect 12032 13572 12036 13628
rect 12036 13572 12092 13628
rect 12092 13572 12096 13628
rect 12032 13568 12096 13572
rect 12112 13628 12176 13632
rect 12112 13572 12116 13628
rect 12116 13572 12172 13628
rect 12172 13572 12176 13628
rect 12112 13568 12176 13572
rect 12192 13628 12256 13632
rect 12192 13572 12196 13628
rect 12196 13572 12252 13628
rect 12252 13572 12256 13628
rect 12192 13568 12256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 21952 13628 22016 13632
rect 21952 13572 21956 13628
rect 21956 13572 22012 13628
rect 22012 13572 22016 13628
rect 21952 13568 22016 13572
rect 22032 13628 22096 13632
rect 22032 13572 22036 13628
rect 22036 13572 22092 13628
rect 22092 13572 22096 13628
rect 22032 13568 22096 13572
rect 22112 13628 22176 13632
rect 22112 13572 22116 13628
rect 22116 13572 22172 13628
rect 22172 13572 22176 13628
rect 22112 13568 22176 13572
rect 22192 13628 22256 13632
rect 22192 13572 22196 13628
rect 22196 13572 22252 13628
rect 22252 13572 22256 13628
rect 22192 13568 22256 13572
rect 26952 13628 27016 13632
rect 26952 13572 26956 13628
rect 26956 13572 27012 13628
rect 27012 13572 27016 13628
rect 26952 13568 27016 13572
rect 27032 13628 27096 13632
rect 27032 13572 27036 13628
rect 27036 13572 27092 13628
rect 27092 13572 27096 13628
rect 27032 13568 27096 13572
rect 27112 13628 27176 13632
rect 27112 13572 27116 13628
rect 27116 13572 27172 13628
rect 27172 13572 27176 13628
rect 27112 13568 27176 13572
rect 27192 13628 27256 13632
rect 27192 13572 27196 13628
rect 27196 13572 27252 13628
rect 27252 13572 27256 13628
rect 27192 13568 27256 13572
rect 31952 13628 32016 13632
rect 31952 13572 31956 13628
rect 31956 13572 32012 13628
rect 32012 13572 32016 13628
rect 31952 13568 32016 13572
rect 32032 13628 32096 13632
rect 32032 13572 32036 13628
rect 32036 13572 32092 13628
rect 32092 13572 32096 13628
rect 32032 13568 32096 13572
rect 32112 13628 32176 13632
rect 32112 13572 32116 13628
rect 32116 13572 32172 13628
rect 32172 13572 32176 13628
rect 32112 13568 32176 13572
rect 32192 13628 32256 13632
rect 32192 13572 32196 13628
rect 32196 13572 32252 13628
rect 32252 13572 32256 13628
rect 32192 13568 32256 13572
rect 36952 13628 37016 13632
rect 36952 13572 36956 13628
rect 36956 13572 37012 13628
rect 37012 13572 37016 13628
rect 36952 13568 37016 13572
rect 37032 13628 37096 13632
rect 37032 13572 37036 13628
rect 37036 13572 37092 13628
rect 37092 13572 37096 13628
rect 37032 13568 37096 13572
rect 37112 13628 37176 13632
rect 37112 13572 37116 13628
rect 37116 13572 37172 13628
rect 37172 13572 37176 13628
rect 37112 13568 37176 13572
rect 37192 13628 37256 13632
rect 37192 13572 37196 13628
rect 37196 13572 37252 13628
rect 37252 13572 37256 13628
rect 37192 13568 37256 13572
rect 2612 13084 2676 13088
rect 2612 13028 2616 13084
rect 2616 13028 2672 13084
rect 2672 13028 2676 13084
rect 2612 13024 2676 13028
rect 2692 13084 2756 13088
rect 2692 13028 2696 13084
rect 2696 13028 2752 13084
rect 2752 13028 2756 13084
rect 2692 13024 2756 13028
rect 2772 13084 2836 13088
rect 2772 13028 2776 13084
rect 2776 13028 2832 13084
rect 2832 13028 2836 13084
rect 2772 13024 2836 13028
rect 2852 13084 2916 13088
rect 2852 13028 2856 13084
rect 2856 13028 2912 13084
rect 2912 13028 2916 13084
rect 2852 13024 2916 13028
rect 7612 13084 7676 13088
rect 7612 13028 7616 13084
rect 7616 13028 7672 13084
rect 7672 13028 7676 13084
rect 7612 13024 7676 13028
rect 7692 13084 7756 13088
rect 7692 13028 7696 13084
rect 7696 13028 7752 13084
rect 7752 13028 7756 13084
rect 7692 13024 7756 13028
rect 7772 13084 7836 13088
rect 7772 13028 7776 13084
rect 7776 13028 7832 13084
rect 7832 13028 7836 13084
rect 7772 13024 7836 13028
rect 7852 13084 7916 13088
rect 7852 13028 7856 13084
rect 7856 13028 7912 13084
rect 7912 13028 7916 13084
rect 7852 13024 7916 13028
rect 12612 13084 12676 13088
rect 12612 13028 12616 13084
rect 12616 13028 12672 13084
rect 12672 13028 12676 13084
rect 12612 13024 12676 13028
rect 12692 13084 12756 13088
rect 12692 13028 12696 13084
rect 12696 13028 12752 13084
rect 12752 13028 12756 13084
rect 12692 13024 12756 13028
rect 12772 13084 12836 13088
rect 12772 13028 12776 13084
rect 12776 13028 12832 13084
rect 12832 13028 12836 13084
rect 12772 13024 12836 13028
rect 12852 13084 12916 13088
rect 12852 13028 12856 13084
rect 12856 13028 12912 13084
rect 12912 13028 12916 13084
rect 12852 13024 12916 13028
rect 17612 13084 17676 13088
rect 17612 13028 17616 13084
rect 17616 13028 17672 13084
rect 17672 13028 17676 13084
rect 17612 13024 17676 13028
rect 17692 13084 17756 13088
rect 17692 13028 17696 13084
rect 17696 13028 17752 13084
rect 17752 13028 17756 13084
rect 17692 13024 17756 13028
rect 17772 13084 17836 13088
rect 17772 13028 17776 13084
rect 17776 13028 17832 13084
rect 17832 13028 17836 13084
rect 17772 13024 17836 13028
rect 17852 13084 17916 13088
rect 17852 13028 17856 13084
rect 17856 13028 17912 13084
rect 17912 13028 17916 13084
rect 17852 13024 17916 13028
rect 22612 13084 22676 13088
rect 22612 13028 22616 13084
rect 22616 13028 22672 13084
rect 22672 13028 22676 13084
rect 22612 13024 22676 13028
rect 22692 13084 22756 13088
rect 22692 13028 22696 13084
rect 22696 13028 22752 13084
rect 22752 13028 22756 13084
rect 22692 13024 22756 13028
rect 22772 13084 22836 13088
rect 22772 13028 22776 13084
rect 22776 13028 22832 13084
rect 22832 13028 22836 13084
rect 22772 13024 22836 13028
rect 22852 13084 22916 13088
rect 22852 13028 22856 13084
rect 22856 13028 22912 13084
rect 22912 13028 22916 13084
rect 22852 13024 22916 13028
rect 27612 13084 27676 13088
rect 27612 13028 27616 13084
rect 27616 13028 27672 13084
rect 27672 13028 27676 13084
rect 27612 13024 27676 13028
rect 27692 13084 27756 13088
rect 27692 13028 27696 13084
rect 27696 13028 27752 13084
rect 27752 13028 27756 13084
rect 27692 13024 27756 13028
rect 27772 13084 27836 13088
rect 27772 13028 27776 13084
rect 27776 13028 27832 13084
rect 27832 13028 27836 13084
rect 27772 13024 27836 13028
rect 27852 13084 27916 13088
rect 27852 13028 27856 13084
rect 27856 13028 27912 13084
rect 27912 13028 27916 13084
rect 27852 13024 27916 13028
rect 32612 13084 32676 13088
rect 32612 13028 32616 13084
rect 32616 13028 32672 13084
rect 32672 13028 32676 13084
rect 32612 13024 32676 13028
rect 32692 13084 32756 13088
rect 32692 13028 32696 13084
rect 32696 13028 32752 13084
rect 32752 13028 32756 13084
rect 32692 13024 32756 13028
rect 32772 13084 32836 13088
rect 32772 13028 32776 13084
rect 32776 13028 32832 13084
rect 32832 13028 32836 13084
rect 32772 13024 32836 13028
rect 32852 13084 32916 13088
rect 32852 13028 32856 13084
rect 32856 13028 32912 13084
rect 32912 13028 32916 13084
rect 32852 13024 32916 13028
rect 37612 13084 37676 13088
rect 37612 13028 37616 13084
rect 37616 13028 37672 13084
rect 37672 13028 37676 13084
rect 37612 13024 37676 13028
rect 37692 13084 37756 13088
rect 37692 13028 37696 13084
rect 37696 13028 37752 13084
rect 37752 13028 37756 13084
rect 37692 13024 37756 13028
rect 37772 13084 37836 13088
rect 37772 13028 37776 13084
rect 37776 13028 37832 13084
rect 37832 13028 37836 13084
rect 37772 13024 37836 13028
rect 37852 13084 37916 13088
rect 37852 13028 37856 13084
rect 37856 13028 37912 13084
rect 37912 13028 37916 13084
rect 37852 13024 37916 13028
rect 1952 12540 2016 12544
rect 1952 12484 1956 12540
rect 1956 12484 2012 12540
rect 2012 12484 2016 12540
rect 1952 12480 2016 12484
rect 2032 12540 2096 12544
rect 2032 12484 2036 12540
rect 2036 12484 2092 12540
rect 2092 12484 2096 12540
rect 2032 12480 2096 12484
rect 2112 12540 2176 12544
rect 2112 12484 2116 12540
rect 2116 12484 2172 12540
rect 2172 12484 2176 12540
rect 2112 12480 2176 12484
rect 2192 12540 2256 12544
rect 2192 12484 2196 12540
rect 2196 12484 2252 12540
rect 2252 12484 2256 12540
rect 2192 12480 2256 12484
rect 6952 12540 7016 12544
rect 6952 12484 6956 12540
rect 6956 12484 7012 12540
rect 7012 12484 7016 12540
rect 6952 12480 7016 12484
rect 7032 12540 7096 12544
rect 7032 12484 7036 12540
rect 7036 12484 7092 12540
rect 7092 12484 7096 12540
rect 7032 12480 7096 12484
rect 7112 12540 7176 12544
rect 7112 12484 7116 12540
rect 7116 12484 7172 12540
rect 7172 12484 7176 12540
rect 7112 12480 7176 12484
rect 7192 12540 7256 12544
rect 7192 12484 7196 12540
rect 7196 12484 7252 12540
rect 7252 12484 7256 12540
rect 7192 12480 7256 12484
rect 11952 12540 12016 12544
rect 11952 12484 11956 12540
rect 11956 12484 12012 12540
rect 12012 12484 12016 12540
rect 11952 12480 12016 12484
rect 12032 12540 12096 12544
rect 12032 12484 12036 12540
rect 12036 12484 12092 12540
rect 12092 12484 12096 12540
rect 12032 12480 12096 12484
rect 12112 12540 12176 12544
rect 12112 12484 12116 12540
rect 12116 12484 12172 12540
rect 12172 12484 12176 12540
rect 12112 12480 12176 12484
rect 12192 12540 12256 12544
rect 12192 12484 12196 12540
rect 12196 12484 12252 12540
rect 12252 12484 12256 12540
rect 12192 12480 12256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 21952 12540 22016 12544
rect 21952 12484 21956 12540
rect 21956 12484 22012 12540
rect 22012 12484 22016 12540
rect 21952 12480 22016 12484
rect 22032 12540 22096 12544
rect 22032 12484 22036 12540
rect 22036 12484 22092 12540
rect 22092 12484 22096 12540
rect 22032 12480 22096 12484
rect 22112 12540 22176 12544
rect 22112 12484 22116 12540
rect 22116 12484 22172 12540
rect 22172 12484 22176 12540
rect 22112 12480 22176 12484
rect 22192 12540 22256 12544
rect 22192 12484 22196 12540
rect 22196 12484 22252 12540
rect 22252 12484 22256 12540
rect 22192 12480 22256 12484
rect 26952 12540 27016 12544
rect 26952 12484 26956 12540
rect 26956 12484 27012 12540
rect 27012 12484 27016 12540
rect 26952 12480 27016 12484
rect 27032 12540 27096 12544
rect 27032 12484 27036 12540
rect 27036 12484 27092 12540
rect 27092 12484 27096 12540
rect 27032 12480 27096 12484
rect 27112 12540 27176 12544
rect 27112 12484 27116 12540
rect 27116 12484 27172 12540
rect 27172 12484 27176 12540
rect 27112 12480 27176 12484
rect 27192 12540 27256 12544
rect 27192 12484 27196 12540
rect 27196 12484 27252 12540
rect 27252 12484 27256 12540
rect 27192 12480 27256 12484
rect 31952 12540 32016 12544
rect 31952 12484 31956 12540
rect 31956 12484 32012 12540
rect 32012 12484 32016 12540
rect 31952 12480 32016 12484
rect 32032 12540 32096 12544
rect 32032 12484 32036 12540
rect 32036 12484 32092 12540
rect 32092 12484 32096 12540
rect 32032 12480 32096 12484
rect 32112 12540 32176 12544
rect 32112 12484 32116 12540
rect 32116 12484 32172 12540
rect 32172 12484 32176 12540
rect 32112 12480 32176 12484
rect 32192 12540 32256 12544
rect 32192 12484 32196 12540
rect 32196 12484 32252 12540
rect 32252 12484 32256 12540
rect 32192 12480 32256 12484
rect 36952 12540 37016 12544
rect 36952 12484 36956 12540
rect 36956 12484 37012 12540
rect 37012 12484 37016 12540
rect 36952 12480 37016 12484
rect 37032 12540 37096 12544
rect 37032 12484 37036 12540
rect 37036 12484 37092 12540
rect 37092 12484 37096 12540
rect 37032 12480 37096 12484
rect 37112 12540 37176 12544
rect 37112 12484 37116 12540
rect 37116 12484 37172 12540
rect 37172 12484 37176 12540
rect 37112 12480 37176 12484
rect 37192 12540 37256 12544
rect 37192 12484 37196 12540
rect 37196 12484 37252 12540
rect 37252 12484 37256 12540
rect 37192 12480 37256 12484
rect 2612 11996 2676 12000
rect 2612 11940 2616 11996
rect 2616 11940 2672 11996
rect 2672 11940 2676 11996
rect 2612 11936 2676 11940
rect 2692 11996 2756 12000
rect 2692 11940 2696 11996
rect 2696 11940 2752 11996
rect 2752 11940 2756 11996
rect 2692 11936 2756 11940
rect 2772 11996 2836 12000
rect 2772 11940 2776 11996
rect 2776 11940 2832 11996
rect 2832 11940 2836 11996
rect 2772 11936 2836 11940
rect 2852 11996 2916 12000
rect 2852 11940 2856 11996
rect 2856 11940 2912 11996
rect 2912 11940 2916 11996
rect 2852 11936 2916 11940
rect 7612 11996 7676 12000
rect 7612 11940 7616 11996
rect 7616 11940 7672 11996
rect 7672 11940 7676 11996
rect 7612 11936 7676 11940
rect 7692 11996 7756 12000
rect 7692 11940 7696 11996
rect 7696 11940 7752 11996
rect 7752 11940 7756 11996
rect 7692 11936 7756 11940
rect 7772 11996 7836 12000
rect 7772 11940 7776 11996
rect 7776 11940 7832 11996
rect 7832 11940 7836 11996
rect 7772 11936 7836 11940
rect 7852 11996 7916 12000
rect 7852 11940 7856 11996
rect 7856 11940 7912 11996
rect 7912 11940 7916 11996
rect 7852 11936 7916 11940
rect 12612 11996 12676 12000
rect 12612 11940 12616 11996
rect 12616 11940 12672 11996
rect 12672 11940 12676 11996
rect 12612 11936 12676 11940
rect 12692 11996 12756 12000
rect 12692 11940 12696 11996
rect 12696 11940 12752 11996
rect 12752 11940 12756 11996
rect 12692 11936 12756 11940
rect 12772 11996 12836 12000
rect 12772 11940 12776 11996
rect 12776 11940 12832 11996
rect 12832 11940 12836 11996
rect 12772 11936 12836 11940
rect 12852 11996 12916 12000
rect 12852 11940 12856 11996
rect 12856 11940 12912 11996
rect 12912 11940 12916 11996
rect 12852 11936 12916 11940
rect 17612 11996 17676 12000
rect 17612 11940 17616 11996
rect 17616 11940 17672 11996
rect 17672 11940 17676 11996
rect 17612 11936 17676 11940
rect 17692 11996 17756 12000
rect 17692 11940 17696 11996
rect 17696 11940 17752 11996
rect 17752 11940 17756 11996
rect 17692 11936 17756 11940
rect 17772 11996 17836 12000
rect 17772 11940 17776 11996
rect 17776 11940 17832 11996
rect 17832 11940 17836 11996
rect 17772 11936 17836 11940
rect 17852 11996 17916 12000
rect 17852 11940 17856 11996
rect 17856 11940 17912 11996
rect 17912 11940 17916 11996
rect 17852 11936 17916 11940
rect 22612 11996 22676 12000
rect 22612 11940 22616 11996
rect 22616 11940 22672 11996
rect 22672 11940 22676 11996
rect 22612 11936 22676 11940
rect 22692 11996 22756 12000
rect 22692 11940 22696 11996
rect 22696 11940 22752 11996
rect 22752 11940 22756 11996
rect 22692 11936 22756 11940
rect 22772 11996 22836 12000
rect 22772 11940 22776 11996
rect 22776 11940 22832 11996
rect 22832 11940 22836 11996
rect 22772 11936 22836 11940
rect 22852 11996 22916 12000
rect 22852 11940 22856 11996
rect 22856 11940 22912 11996
rect 22912 11940 22916 11996
rect 22852 11936 22916 11940
rect 27612 11996 27676 12000
rect 27612 11940 27616 11996
rect 27616 11940 27672 11996
rect 27672 11940 27676 11996
rect 27612 11936 27676 11940
rect 27692 11996 27756 12000
rect 27692 11940 27696 11996
rect 27696 11940 27752 11996
rect 27752 11940 27756 11996
rect 27692 11936 27756 11940
rect 27772 11996 27836 12000
rect 27772 11940 27776 11996
rect 27776 11940 27832 11996
rect 27832 11940 27836 11996
rect 27772 11936 27836 11940
rect 27852 11996 27916 12000
rect 27852 11940 27856 11996
rect 27856 11940 27912 11996
rect 27912 11940 27916 11996
rect 27852 11936 27916 11940
rect 32612 11996 32676 12000
rect 32612 11940 32616 11996
rect 32616 11940 32672 11996
rect 32672 11940 32676 11996
rect 32612 11936 32676 11940
rect 32692 11996 32756 12000
rect 32692 11940 32696 11996
rect 32696 11940 32752 11996
rect 32752 11940 32756 11996
rect 32692 11936 32756 11940
rect 32772 11996 32836 12000
rect 32772 11940 32776 11996
rect 32776 11940 32832 11996
rect 32832 11940 32836 11996
rect 32772 11936 32836 11940
rect 32852 11996 32916 12000
rect 32852 11940 32856 11996
rect 32856 11940 32912 11996
rect 32912 11940 32916 11996
rect 32852 11936 32916 11940
rect 37612 11996 37676 12000
rect 37612 11940 37616 11996
rect 37616 11940 37672 11996
rect 37672 11940 37676 11996
rect 37612 11936 37676 11940
rect 37692 11996 37756 12000
rect 37692 11940 37696 11996
rect 37696 11940 37752 11996
rect 37752 11940 37756 11996
rect 37692 11936 37756 11940
rect 37772 11996 37836 12000
rect 37772 11940 37776 11996
rect 37776 11940 37832 11996
rect 37832 11940 37836 11996
rect 37772 11936 37836 11940
rect 37852 11996 37916 12000
rect 37852 11940 37856 11996
rect 37856 11940 37912 11996
rect 37912 11940 37916 11996
rect 37852 11936 37916 11940
rect 1952 11452 2016 11456
rect 1952 11396 1956 11452
rect 1956 11396 2012 11452
rect 2012 11396 2016 11452
rect 1952 11392 2016 11396
rect 2032 11452 2096 11456
rect 2032 11396 2036 11452
rect 2036 11396 2092 11452
rect 2092 11396 2096 11452
rect 2032 11392 2096 11396
rect 2112 11452 2176 11456
rect 2112 11396 2116 11452
rect 2116 11396 2172 11452
rect 2172 11396 2176 11452
rect 2112 11392 2176 11396
rect 2192 11452 2256 11456
rect 2192 11396 2196 11452
rect 2196 11396 2252 11452
rect 2252 11396 2256 11452
rect 2192 11392 2256 11396
rect 6952 11452 7016 11456
rect 6952 11396 6956 11452
rect 6956 11396 7012 11452
rect 7012 11396 7016 11452
rect 6952 11392 7016 11396
rect 7032 11452 7096 11456
rect 7032 11396 7036 11452
rect 7036 11396 7092 11452
rect 7092 11396 7096 11452
rect 7032 11392 7096 11396
rect 7112 11452 7176 11456
rect 7112 11396 7116 11452
rect 7116 11396 7172 11452
rect 7172 11396 7176 11452
rect 7112 11392 7176 11396
rect 7192 11452 7256 11456
rect 7192 11396 7196 11452
rect 7196 11396 7252 11452
rect 7252 11396 7256 11452
rect 7192 11392 7256 11396
rect 11952 11452 12016 11456
rect 11952 11396 11956 11452
rect 11956 11396 12012 11452
rect 12012 11396 12016 11452
rect 11952 11392 12016 11396
rect 12032 11452 12096 11456
rect 12032 11396 12036 11452
rect 12036 11396 12092 11452
rect 12092 11396 12096 11452
rect 12032 11392 12096 11396
rect 12112 11452 12176 11456
rect 12112 11396 12116 11452
rect 12116 11396 12172 11452
rect 12172 11396 12176 11452
rect 12112 11392 12176 11396
rect 12192 11452 12256 11456
rect 12192 11396 12196 11452
rect 12196 11396 12252 11452
rect 12252 11396 12256 11452
rect 12192 11392 12256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 21952 11452 22016 11456
rect 21952 11396 21956 11452
rect 21956 11396 22012 11452
rect 22012 11396 22016 11452
rect 21952 11392 22016 11396
rect 22032 11452 22096 11456
rect 22032 11396 22036 11452
rect 22036 11396 22092 11452
rect 22092 11396 22096 11452
rect 22032 11392 22096 11396
rect 22112 11452 22176 11456
rect 22112 11396 22116 11452
rect 22116 11396 22172 11452
rect 22172 11396 22176 11452
rect 22112 11392 22176 11396
rect 22192 11452 22256 11456
rect 22192 11396 22196 11452
rect 22196 11396 22252 11452
rect 22252 11396 22256 11452
rect 22192 11392 22256 11396
rect 26952 11452 27016 11456
rect 26952 11396 26956 11452
rect 26956 11396 27012 11452
rect 27012 11396 27016 11452
rect 26952 11392 27016 11396
rect 27032 11452 27096 11456
rect 27032 11396 27036 11452
rect 27036 11396 27092 11452
rect 27092 11396 27096 11452
rect 27032 11392 27096 11396
rect 27112 11452 27176 11456
rect 27112 11396 27116 11452
rect 27116 11396 27172 11452
rect 27172 11396 27176 11452
rect 27112 11392 27176 11396
rect 27192 11452 27256 11456
rect 27192 11396 27196 11452
rect 27196 11396 27252 11452
rect 27252 11396 27256 11452
rect 27192 11392 27256 11396
rect 31952 11452 32016 11456
rect 31952 11396 31956 11452
rect 31956 11396 32012 11452
rect 32012 11396 32016 11452
rect 31952 11392 32016 11396
rect 32032 11452 32096 11456
rect 32032 11396 32036 11452
rect 32036 11396 32092 11452
rect 32092 11396 32096 11452
rect 32032 11392 32096 11396
rect 32112 11452 32176 11456
rect 32112 11396 32116 11452
rect 32116 11396 32172 11452
rect 32172 11396 32176 11452
rect 32112 11392 32176 11396
rect 32192 11452 32256 11456
rect 32192 11396 32196 11452
rect 32196 11396 32252 11452
rect 32252 11396 32256 11452
rect 32192 11392 32256 11396
rect 36952 11452 37016 11456
rect 36952 11396 36956 11452
rect 36956 11396 37012 11452
rect 37012 11396 37016 11452
rect 36952 11392 37016 11396
rect 37032 11452 37096 11456
rect 37032 11396 37036 11452
rect 37036 11396 37092 11452
rect 37092 11396 37096 11452
rect 37032 11392 37096 11396
rect 37112 11452 37176 11456
rect 37112 11396 37116 11452
rect 37116 11396 37172 11452
rect 37172 11396 37176 11452
rect 37112 11392 37176 11396
rect 37192 11452 37256 11456
rect 37192 11396 37196 11452
rect 37196 11396 37252 11452
rect 37252 11396 37256 11452
rect 37192 11392 37256 11396
rect 2612 10908 2676 10912
rect 2612 10852 2616 10908
rect 2616 10852 2672 10908
rect 2672 10852 2676 10908
rect 2612 10848 2676 10852
rect 2692 10908 2756 10912
rect 2692 10852 2696 10908
rect 2696 10852 2752 10908
rect 2752 10852 2756 10908
rect 2692 10848 2756 10852
rect 2772 10908 2836 10912
rect 2772 10852 2776 10908
rect 2776 10852 2832 10908
rect 2832 10852 2836 10908
rect 2772 10848 2836 10852
rect 2852 10908 2916 10912
rect 2852 10852 2856 10908
rect 2856 10852 2912 10908
rect 2912 10852 2916 10908
rect 2852 10848 2916 10852
rect 7612 10908 7676 10912
rect 7612 10852 7616 10908
rect 7616 10852 7672 10908
rect 7672 10852 7676 10908
rect 7612 10848 7676 10852
rect 7692 10908 7756 10912
rect 7692 10852 7696 10908
rect 7696 10852 7752 10908
rect 7752 10852 7756 10908
rect 7692 10848 7756 10852
rect 7772 10908 7836 10912
rect 7772 10852 7776 10908
rect 7776 10852 7832 10908
rect 7832 10852 7836 10908
rect 7772 10848 7836 10852
rect 7852 10908 7916 10912
rect 7852 10852 7856 10908
rect 7856 10852 7912 10908
rect 7912 10852 7916 10908
rect 7852 10848 7916 10852
rect 12612 10908 12676 10912
rect 12612 10852 12616 10908
rect 12616 10852 12672 10908
rect 12672 10852 12676 10908
rect 12612 10848 12676 10852
rect 12692 10908 12756 10912
rect 12692 10852 12696 10908
rect 12696 10852 12752 10908
rect 12752 10852 12756 10908
rect 12692 10848 12756 10852
rect 12772 10908 12836 10912
rect 12772 10852 12776 10908
rect 12776 10852 12832 10908
rect 12832 10852 12836 10908
rect 12772 10848 12836 10852
rect 12852 10908 12916 10912
rect 12852 10852 12856 10908
rect 12856 10852 12912 10908
rect 12912 10852 12916 10908
rect 12852 10848 12916 10852
rect 17612 10908 17676 10912
rect 17612 10852 17616 10908
rect 17616 10852 17672 10908
rect 17672 10852 17676 10908
rect 17612 10848 17676 10852
rect 17692 10908 17756 10912
rect 17692 10852 17696 10908
rect 17696 10852 17752 10908
rect 17752 10852 17756 10908
rect 17692 10848 17756 10852
rect 17772 10908 17836 10912
rect 17772 10852 17776 10908
rect 17776 10852 17832 10908
rect 17832 10852 17836 10908
rect 17772 10848 17836 10852
rect 17852 10908 17916 10912
rect 17852 10852 17856 10908
rect 17856 10852 17912 10908
rect 17912 10852 17916 10908
rect 17852 10848 17916 10852
rect 22612 10908 22676 10912
rect 22612 10852 22616 10908
rect 22616 10852 22672 10908
rect 22672 10852 22676 10908
rect 22612 10848 22676 10852
rect 22692 10908 22756 10912
rect 22692 10852 22696 10908
rect 22696 10852 22752 10908
rect 22752 10852 22756 10908
rect 22692 10848 22756 10852
rect 22772 10908 22836 10912
rect 22772 10852 22776 10908
rect 22776 10852 22832 10908
rect 22832 10852 22836 10908
rect 22772 10848 22836 10852
rect 22852 10908 22916 10912
rect 22852 10852 22856 10908
rect 22856 10852 22912 10908
rect 22912 10852 22916 10908
rect 22852 10848 22916 10852
rect 27612 10908 27676 10912
rect 27612 10852 27616 10908
rect 27616 10852 27672 10908
rect 27672 10852 27676 10908
rect 27612 10848 27676 10852
rect 27692 10908 27756 10912
rect 27692 10852 27696 10908
rect 27696 10852 27752 10908
rect 27752 10852 27756 10908
rect 27692 10848 27756 10852
rect 27772 10908 27836 10912
rect 27772 10852 27776 10908
rect 27776 10852 27832 10908
rect 27832 10852 27836 10908
rect 27772 10848 27836 10852
rect 27852 10908 27916 10912
rect 27852 10852 27856 10908
rect 27856 10852 27912 10908
rect 27912 10852 27916 10908
rect 27852 10848 27916 10852
rect 32612 10908 32676 10912
rect 32612 10852 32616 10908
rect 32616 10852 32672 10908
rect 32672 10852 32676 10908
rect 32612 10848 32676 10852
rect 32692 10908 32756 10912
rect 32692 10852 32696 10908
rect 32696 10852 32752 10908
rect 32752 10852 32756 10908
rect 32692 10848 32756 10852
rect 32772 10908 32836 10912
rect 32772 10852 32776 10908
rect 32776 10852 32832 10908
rect 32832 10852 32836 10908
rect 32772 10848 32836 10852
rect 32852 10908 32916 10912
rect 32852 10852 32856 10908
rect 32856 10852 32912 10908
rect 32912 10852 32916 10908
rect 32852 10848 32916 10852
rect 37612 10908 37676 10912
rect 37612 10852 37616 10908
rect 37616 10852 37672 10908
rect 37672 10852 37676 10908
rect 37612 10848 37676 10852
rect 37692 10908 37756 10912
rect 37692 10852 37696 10908
rect 37696 10852 37752 10908
rect 37752 10852 37756 10908
rect 37692 10848 37756 10852
rect 37772 10908 37836 10912
rect 37772 10852 37776 10908
rect 37776 10852 37832 10908
rect 37832 10852 37836 10908
rect 37772 10848 37836 10852
rect 37852 10908 37916 10912
rect 37852 10852 37856 10908
rect 37856 10852 37912 10908
rect 37912 10852 37916 10908
rect 37852 10848 37916 10852
rect 1952 10364 2016 10368
rect 1952 10308 1956 10364
rect 1956 10308 2012 10364
rect 2012 10308 2016 10364
rect 1952 10304 2016 10308
rect 2032 10364 2096 10368
rect 2032 10308 2036 10364
rect 2036 10308 2092 10364
rect 2092 10308 2096 10364
rect 2032 10304 2096 10308
rect 2112 10364 2176 10368
rect 2112 10308 2116 10364
rect 2116 10308 2172 10364
rect 2172 10308 2176 10364
rect 2112 10304 2176 10308
rect 2192 10364 2256 10368
rect 2192 10308 2196 10364
rect 2196 10308 2252 10364
rect 2252 10308 2256 10364
rect 2192 10304 2256 10308
rect 6952 10364 7016 10368
rect 6952 10308 6956 10364
rect 6956 10308 7012 10364
rect 7012 10308 7016 10364
rect 6952 10304 7016 10308
rect 7032 10364 7096 10368
rect 7032 10308 7036 10364
rect 7036 10308 7092 10364
rect 7092 10308 7096 10364
rect 7032 10304 7096 10308
rect 7112 10364 7176 10368
rect 7112 10308 7116 10364
rect 7116 10308 7172 10364
rect 7172 10308 7176 10364
rect 7112 10304 7176 10308
rect 7192 10364 7256 10368
rect 7192 10308 7196 10364
rect 7196 10308 7252 10364
rect 7252 10308 7256 10364
rect 7192 10304 7256 10308
rect 11952 10364 12016 10368
rect 11952 10308 11956 10364
rect 11956 10308 12012 10364
rect 12012 10308 12016 10364
rect 11952 10304 12016 10308
rect 12032 10364 12096 10368
rect 12032 10308 12036 10364
rect 12036 10308 12092 10364
rect 12092 10308 12096 10364
rect 12032 10304 12096 10308
rect 12112 10364 12176 10368
rect 12112 10308 12116 10364
rect 12116 10308 12172 10364
rect 12172 10308 12176 10364
rect 12112 10304 12176 10308
rect 12192 10364 12256 10368
rect 12192 10308 12196 10364
rect 12196 10308 12252 10364
rect 12252 10308 12256 10364
rect 12192 10304 12256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 21952 10364 22016 10368
rect 21952 10308 21956 10364
rect 21956 10308 22012 10364
rect 22012 10308 22016 10364
rect 21952 10304 22016 10308
rect 22032 10364 22096 10368
rect 22032 10308 22036 10364
rect 22036 10308 22092 10364
rect 22092 10308 22096 10364
rect 22032 10304 22096 10308
rect 22112 10364 22176 10368
rect 22112 10308 22116 10364
rect 22116 10308 22172 10364
rect 22172 10308 22176 10364
rect 22112 10304 22176 10308
rect 22192 10364 22256 10368
rect 22192 10308 22196 10364
rect 22196 10308 22252 10364
rect 22252 10308 22256 10364
rect 22192 10304 22256 10308
rect 26952 10364 27016 10368
rect 26952 10308 26956 10364
rect 26956 10308 27012 10364
rect 27012 10308 27016 10364
rect 26952 10304 27016 10308
rect 27032 10364 27096 10368
rect 27032 10308 27036 10364
rect 27036 10308 27092 10364
rect 27092 10308 27096 10364
rect 27032 10304 27096 10308
rect 27112 10364 27176 10368
rect 27112 10308 27116 10364
rect 27116 10308 27172 10364
rect 27172 10308 27176 10364
rect 27112 10304 27176 10308
rect 27192 10364 27256 10368
rect 27192 10308 27196 10364
rect 27196 10308 27252 10364
rect 27252 10308 27256 10364
rect 27192 10304 27256 10308
rect 31952 10364 32016 10368
rect 31952 10308 31956 10364
rect 31956 10308 32012 10364
rect 32012 10308 32016 10364
rect 31952 10304 32016 10308
rect 32032 10364 32096 10368
rect 32032 10308 32036 10364
rect 32036 10308 32092 10364
rect 32092 10308 32096 10364
rect 32032 10304 32096 10308
rect 32112 10364 32176 10368
rect 32112 10308 32116 10364
rect 32116 10308 32172 10364
rect 32172 10308 32176 10364
rect 32112 10304 32176 10308
rect 32192 10364 32256 10368
rect 32192 10308 32196 10364
rect 32196 10308 32252 10364
rect 32252 10308 32256 10364
rect 32192 10304 32256 10308
rect 36952 10364 37016 10368
rect 36952 10308 36956 10364
rect 36956 10308 37012 10364
rect 37012 10308 37016 10364
rect 36952 10304 37016 10308
rect 37032 10364 37096 10368
rect 37032 10308 37036 10364
rect 37036 10308 37092 10364
rect 37092 10308 37096 10364
rect 37032 10304 37096 10308
rect 37112 10364 37176 10368
rect 37112 10308 37116 10364
rect 37116 10308 37172 10364
rect 37172 10308 37176 10364
rect 37112 10304 37176 10308
rect 37192 10364 37256 10368
rect 37192 10308 37196 10364
rect 37196 10308 37252 10364
rect 37252 10308 37256 10364
rect 37192 10304 37256 10308
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 7612 9820 7676 9824
rect 7612 9764 7616 9820
rect 7616 9764 7672 9820
rect 7672 9764 7676 9820
rect 7612 9760 7676 9764
rect 7692 9820 7756 9824
rect 7692 9764 7696 9820
rect 7696 9764 7752 9820
rect 7752 9764 7756 9820
rect 7692 9760 7756 9764
rect 7772 9820 7836 9824
rect 7772 9764 7776 9820
rect 7776 9764 7832 9820
rect 7832 9764 7836 9820
rect 7772 9760 7836 9764
rect 7852 9820 7916 9824
rect 7852 9764 7856 9820
rect 7856 9764 7912 9820
rect 7912 9764 7916 9820
rect 7852 9760 7916 9764
rect 12612 9820 12676 9824
rect 12612 9764 12616 9820
rect 12616 9764 12672 9820
rect 12672 9764 12676 9820
rect 12612 9760 12676 9764
rect 12692 9820 12756 9824
rect 12692 9764 12696 9820
rect 12696 9764 12752 9820
rect 12752 9764 12756 9820
rect 12692 9760 12756 9764
rect 12772 9820 12836 9824
rect 12772 9764 12776 9820
rect 12776 9764 12832 9820
rect 12832 9764 12836 9820
rect 12772 9760 12836 9764
rect 12852 9820 12916 9824
rect 12852 9764 12856 9820
rect 12856 9764 12912 9820
rect 12912 9764 12916 9820
rect 12852 9760 12916 9764
rect 17612 9820 17676 9824
rect 17612 9764 17616 9820
rect 17616 9764 17672 9820
rect 17672 9764 17676 9820
rect 17612 9760 17676 9764
rect 17692 9820 17756 9824
rect 17692 9764 17696 9820
rect 17696 9764 17752 9820
rect 17752 9764 17756 9820
rect 17692 9760 17756 9764
rect 17772 9820 17836 9824
rect 17772 9764 17776 9820
rect 17776 9764 17832 9820
rect 17832 9764 17836 9820
rect 17772 9760 17836 9764
rect 17852 9820 17916 9824
rect 17852 9764 17856 9820
rect 17856 9764 17912 9820
rect 17912 9764 17916 9820
rect 17852 9760 17916 9764
rect 22612 9820 22676 9824
rect 22612 9764 22616 9820
rect 22616 9764 22672 9820
rect 22672 9764 22676 9820
rect 22612 9760 22676 9764
rect 22692 9820 22756 9824
rect 22692 9764 22696 9820
rect 22696 9764 22752 9820
rect 22752 9764 22756 9820
rect 22692 9760 22756 9764
rect 22772 9820 22836 9824
rect 22772 9764 22776 9820
rect 22776 9764 22832 9820
rect 22832 9764 22836 9820
rect 22772 9760 22836 9764
rect 22852 9820 22916 9824
rect 22852 9764 22856 9820
rect 22856 9764 22912 9820
rect 22912 9764 22916 9820
rect 22852 9760 22916 9764
rect 27612 9820 27676 9824
rect 27612 9764 27616 9820
rect 27616 9764 27672 9820
rect 27672 9764 27676 9820
rect 27612 9760 27676 9764
rect 27692 9820 27756 9824
rect 27692 9764 27696 9820
rect 27696 9764 27752 9820
rect 27752 9764 27756 9820
rect 27692 9760 27756 9764
rect 27772 9820 27836 9824
rect 27772 9764 27776 9820
rect 27776 9764 27832 9820
rect 27832 9764 27836 9820
rect 27772 9760 27836 9764
rect 27852 9820 27916 9824
rect 27852 9764 27856 9820
rect 27856 9764 27912 9820
rect 27912 9764 27916 9820
rect 27852 9760 27916 9764
rect 32612 9820 32676 9824
rect 32612 9764 32616 9820
rect 32616 9764 32672 9820
rect 32672 9764 32676 9820
rect 32612 9760 32676 9764
rect 32692 9820 32756 9824
rect 32692 9764 32696 9820
rect 32696 9764 32752 9820
rect 32752 9764 32756 9820
rect 32692 9760 32756 9764
rect 32772 9820 32836 9824
rect 32772 9764 32776 9820
rect 32776 9764 32832 9820
rect 32832 9764 32836 9820
rect 32772 9760 32836 9764
rect 32852 9820 32916 9824
rect 32852 9764 32856 9820
rect 32856 9764 32912 9820
rect 32912 9764 32916 9820
rect 32852 9760 32916 9764
rect 37612 9820 37676 9824
rect 37612 9764 37616 9820
rect 37616 9764 37672 9820
rect 37672 9764 37676 9820
rect 37612 9760 37676 9764
rect 37692 9820 37756 9824
rect 37692 9764 37696 9820
rect 37696 9764 37752 9820
rect 37752 9764 37756 9820
rect 37692 9760 37756 9764
rect 37772 9820 37836 9824
rect 37772 9764 37776 9820
rect 37776 9764 37832 9820
rect 37832 9764 37836 9820
rect 37772 9760 37836 9764
rect 37852 9820 37916 9824
rect 37852 9764 37856 9820
rect 37856 9764 37912 9820
rect 37912 9764 37916 9820
rect 37852 9760 37916 9764
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 6952 9276 7016 9280
rect 6952 9220 6956 9276
rect 6956 9220 7012 9276
rect 7012 9220 7016 9276
rect 6952 9216 7016 9220
rect 7032 9276 7096 9280
rect 7032 9220 7036 9276
rect 7036 9220 7092 9276
rect 7092 9220 7096 9276
rect 7032 9216 7096 9220
rect 7112 9276 7176 9280
rect 7112 9220 7116 9276
rect 7116 9220 7172 9276
rect 7172 9220 7176 9276
rect 7112 9216 7176 9220
rect 7192 9276 7256 9280
rect 7192 9220 7196 9276
rect 7196 9220 7252 9276
rect 7252 9220 7256 9276
rect 7192 9216 7256 9220
rect 11952 9276 12016 9280
rect 11952 9220 11956 9276
rect 11956 9220 12012 9276
rect 12012 9220 12016 9276
rect 11952 9216 12016 9220
rect 12032 9276 12096 9280
rect 12032 9220 12036 9276
rect 12036 9220 12092 9276
rect 12092 9220 12096 9276
rect 12032 9216 12096 9220
rect 12112 9276 12176 9280
rect 12112 9220 12116 9276
rect 12116 9220 12172 9276
rect 12172 9220 12176 9276
rect 12112 9216 12176 9220
rect 12192 9276 12256 9280
rect 12192 9220 12196 9276
rect 12196 9220 12252 9276
rect 12252 9220 12256 9276
rect 12192 9216 12256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 21952 9276 22016 9280
rect 21952 9220 21956 9276
rect 21956 9220 22012 9276
rect 22012 9220 22016 9276
rect 21952 9216 22016 9220
rect 22032 9276 22096 9280
rect 22032 9220 22036 9276
rect 22036 9220 22092 9276
rect 22092 9220 22096 9276
rect 22032 9216 22096 9220
rect 22112 9276 22176 9280
rect 22112 9220 22116 9276
rect 22116 9220 22172 9276
rect 22172 9220 22176 9276
rect 22112 9216 22176 9220
rect 22192 9276 22256 9280
rect 22192 9220 22196 9276
rect 22196 9220 22252 9276
rect 22252 9220 22256 9276
rect 22192 9216 22256 9220
rect 26952 9276 27016 9280
rect 26952 9220 26956 9276
rect 26956 9220 27012 9276
rect 27012 9220 27016 9276
rect 26952 9216 27016 9220
rect 27032 9276 27096 9280
rect 27032 9220 27036 9276
rect 27036 9220 27092 9276
rect 27092 9220 27096 9276
rect 27032 9216 27096 9220
rect 27112 9276 27176 9280
rect 27112 9220 27116 9276
rect 27116 9220 27172 9276
rect 27172 9220 27176 9276
rect 27112 9216 27176 9220
rect 27192 9276 27256 9280
rect 27192 9220 27196 9276
rect 27196 9220 27252 9276
rect 27252 9220 27256 9276
rect 27192 9216 27256 9220
rect 31952 9276 32016 9280
rect 31952 9220 31956 9276
rect 31956 9220 32012 9276
rect 32012 9220 32016 9276
rect 31952 9216 32016 9220
rect 32032 9276 32096 9280
rect 32032 9220 32036 9276
rect 32036 9220 32092 9276
rect 32092 9220 32096 9276
rect 32032 9216 32096 9220
rect 32112 9276 32176 9280
rect 32112 9220 32116 9276
rect 32116 9220 32172 9276
rect 32172 9220 32176 9276
rect 32112 9216 32176 9220
rect 32192 9276 32256 9280
rect 32192 9220 32196 9276
rect 32196 9220 32252 9276
rect 32252 9220 32256 9276
rect 32192 9216 32256 9220
rect 36952 9276 37016 9280
rect 36952 9220 36956 9276
rect 36956 9220 37012 9276
rect 37012 9220 37016 9276
rect 36952 9216 37016 9220
rect 37032 9276 37096 9280
rect 37032 9220 37036 9276
rect 37036 9220 37092 9276
rect 37092 9220 37096 9276
rect 37032 9216 37096 9220
rect 37112 9276 37176 9280
rect 37112 9220 37116 9276
rect 37116 9220 37172 9276
rect 37172 9220 37176 9276
rect 37112 9216 37176 9220
rect 37192 9276 37256 9280
rect 37192 9220 37196 9276
rect 37196 9220 37252 9276
rect 37252 9220 37256 9276
rect 37192 9216 37256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 7612 8732 7676 8736
rect 7612 8676 7616 8732
rect 7616 8676 7672 8732
rect 7672 8676 7676 8732
rect 7612 8672 7676 8676
rect 7692 8732 7756 8736
rect 7692 8676 7696 8732
rect 7696 8676 7752 8732
rect 7752 8676 7756 8732
rect 7692 8672 7756 8676
rect 7772 8732 7836 8736
rect 7772 8676 7776 8732
rect 7776 8676 7832 8732
rect 7832 8676 7836 8732
rect 7772 8672 7836 8676
rect 7852 8732 7916 8736
rect 7852 8676 7856 8732
rect 7856 8676 7912 8732
rect 7912 8676 7916 8732
rect 7852 8672 7916 8676
rect 12612 8732 12676 8736
rect 12612 8676 12616 8732
rect 12616 8676 12672 8732
rect 12672 8676 12676 8732
rect 12612 8672 12676 8676
rect 12692 8732 12756 8736
rect 12692 8676 12696 8732
rect 12696 8676 12752 8732
rect 12752 8676 12756 8732
rect 12692 8672 12756 8676
rect 12772 8732 12836 8736
rect 12772 8676 12776 8732
rect 12776 8676 12832 8732
rect 12832 8676 12836 8732
rect 12772 8672 12836 8676
rect 12852 8732 12916 8736
rect 12852 8676 12856 8732
rect 12856 8676 12912 8732
rect 12912 8676 12916 8732
rect 12852 8672 12916 8676
rect 17612 8732 17676 8736
rect 17612 8676 17616 8732
rect 17616 8676 17672 8732
rect 17672 8676 17676 8732
rect 17612 8672 17676 8676
rect 17692 8732 17756 8736
rect 17692 8676 17696 8732
rect 17696 8676 17752 8732
rect 17752 8676 17756 8732
rect 17692 8672 17756 8676
rect 17772 8732 17836 8736
rect 17772 8676 17776 8732
rect 17776 8676 17832 8732
rect 17832 8676 17836 8732
rect 17772 8672 17836 8676
rect 17852 8732 17916 8736
rect 17852 8676 17856 8732
rect 17856 8676 17912 8732
rect 17912 8676 17916 8732
rect 17852 8672 17916 8676
rect 22612 8732 22676 8736
rect 22612 8676 22616 8732
rect 22616 8676 22672 8732
rect 22672 8676 22676 8732
rect 22612 8672 22676 8676
rect 22692 8732 22756 8736
rect 22692 8676 22696 8732
rect 22696 8676 22752 8732
rect 22752 8676 22756 8732
rect 22692 8672 22756 8676
rect 22772 8732 22836 8736
rect 22772 8676 22776 8732
rect 22776 8676 22832 8732
rect 22832 8676 22836 8732
rect 22772 8672 22836 8676
rect 22852 8732 22916 8736
rect 22852 8676 22856 8732
rect 22856 8676 22912 8732
rect 22912 8676 22916 8732
rect 22852 8672 22916 8676
rect 27612 8732 27676 8736
rect 27612 8676 27616 8732
rect 27616 8676 27672 8732
rect 27672 8676 27676 8732
rect 27612 8672 27676 8676
rect 27692 8732 27756 8736
rect 27692 8676 27696 8732
rect 27696 8676 27752 8732
rect 27752 8676 27756 8732
rect 27692 8672 27756 8676
rect 27772 8732 27836 8736
rect 27772 8676 27776 8732
rect 27776 8676 27832 8732
rect 27832 8676 27836 8732
rect 27772 8672 27836 8676
rect 27852 8732 27916 8736
rect 27852 8676 27856 8732
rect 27856 8676 27912 8732
rect 27912 8676 27916 8732
rect 27852 8672 27916 8676
rect 32612 8732 32676 8736
rect 32612 8676 32616 8732
rect 32616 8676 32672 8732
rect 32672 8676 32676 8732
rect 32612 8672 32676 8676
rect 32692 8732 32756 8736
rect 32692 8676 32696 8732
rect 32696 8676 32752 8732
rect 32752 8676 32756 8732
rect 32692 8672 32756 8676
rect 32772 8732 32836 8736
rect 32772 8676 32776 8732
rect 32776 8676 32832 8732
rect 32832 8676 32836 8732
rect 32772 8672 32836 8676
rect 32852 8732 32916 8736
rect 32852 8676 32856 8732
rect 32856 8676 32912 8732
rect 32912 8676 32916 8732
rect 32852 8672 32916 8676
rect 37612 8732 37676 8736
rect 37612 8676 37616 8732
rect 37616 8676 37672 8732
rect 37672 8676 37676 8732
rect 37612 8672 37676 8676
rect 37692 8732 37756 8736
rect 37692 8676 37696 8732
rect 37696 8676 37752 8732
rect 37752 8676 37756 8732
rect 37692 8672 37756 8676
rect 37772 8732 37836 8736
rect 37772 8676 37776 8732
rect 37776 8676 37832 8732
rect 37832 8676 37836 8732
rect 37772 8672 37836 8676
rect 37852 8732 37916 8736
rect 37852 8676 37856 8732
rect 37856 8676 37912 8732
rect 37912 8676 37916 8732
rect 37852 8672 37916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 6952 8188 7016 8192
rect 6952 8132 6956 8188
rect 6956 8132 7012 8188
rect 7012 8132 7016 8188
rect 6952 8128 7016 8132
rect 7032 8188 7096 8192
rect 7032 8132 7036 8188
rect 7036 8132 7092 8188
rect 7092 8132 7096 8188
rect 7032 8128 7096 8132
rect 7112 8188 7176 8192
rect 7112 8132 7116 8188
rect 7116 8132 7172 8188
rect 7172 8132 7176 8188
rect 7112 8128 7176 8132
rect 7192 8188 7256 8192
rect 7192 8132 7196 8188
rect 7196 8132 7252 8188
rect 7252 8132 7256 8188
rect 7192 8128 7256 8132
rect 11952 8188 12016 8192
rect 11952 8132 11956 8188
rect 11956 8132 12012 8188
rect 12012 8132 12016 8188
rect 11952 8128 12016 8132
rect 12032 8188 12096 8192
rect 12032 8132 12036 8188
rect 12036 8132 12092 8188
rect 12092 8132 12096 8188
rect 12032 8128 12096 8132
rect 12112 8188 12176 8192
rect 12112 8132 12116 8188
rect 12116 8132 12172 8188
rect 12172 8132 12176 8188
rect 12112 8128 12176 8132
rect 12192 8188 12256 8192
rect 12192 8132 12196 8188
rect 12196 8132 12252 8188
rect 12252 8132 12256 8188
rect 12192 8128 12256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 21952 8188 22016 8192
rect 21952 8132 21956 8188
rect 21956 8132 22012 8188
rect 22012 8132 22016 8188
rect 21952 8128 22016 8132
rect 22032 8188 22096 8192
rect 22032 8132 22036 8188
rect 22036 8132 22092 8188
rect 22092 8132 22096 8188
rect 22032 8128 22096 8132
rect 22112 8188 22176 8192
rect 22112 8132 22116 8188
rect 22116 8132 22172 8188
rect 22172 8132 22176 8188
rect 22112 8128 22176 8132
rect 22192 8188 22256 8192
rect 22192 8132 22196 8188
rect 22196 8132 22252 8188
rect 22252 8132 22256 8188
rect 22192 8128 22256 8132
rect 26952 8188 27016 8192
rect 26952 8132 26956 8188
rect 26956 8132 27012 8188
rect 27012 8132 27016 8188
rect 26952 8128 27016 8132
rect 27032 8188 27096 8192
rect 27032 8132 27036 8188
rect 27036 8132 27092 8188
rect 27092 8132 27096 8188
rect 27032 8128 27096 8132
rect 27112 8188 27176 8192
rect 27112 8132 27116 8188
rect 27116 8132 27172 8188
rect 27172 8132 27176 8188
rect 27112 8128 27176 8132
rect 27192 8188 27256 8192
rect 27192 8132 27196 8188
rect 27196 8132 27252 8188
rect 27252 8132 27256 8188
rect 27192 8128 27256 8132
rect 31952 8188 32016 8192
rect 31952 8132 31956 8188
rect 31956 8132 32012 8188
rect 32012 8132 32016 8188
rect 31952 8128 32016 8132
rect 32032 8188 32096 8192
rect 32032 8132 32036 8188
rect 32036 8132 32092 8188
rect 32092 8132 32096 8188
rect 32032 8128 32096 8132
rect 32112 8188 32176 8192
rect 32112 8132 32116 8188
rect 32116 8132 32172 8188
rect 32172 8132 32176 8188
rect 32112 8128 32176 8132
rect 32192 8188 32256 8192
rect 32192 8132 32196 8188
rect 32196 8132 32252 8188
rect 32252 8132 32256 8188
rect 32192 8128 32256 8132
rect 36952 8188 37016 8192
rect 36952 8132 36956 8188
rect 36956 8132 37012 8188
rect 37012 8132 37016 8188
rect 36952 8128 37016 8132
rect 37032 8188 37096 8192
rect 37032 8132 37036 8188
rect 37036 8132 37092 8188
rect 37092 8132 37096 8188
rect 37032 8128 37096 8132
rect 37112 8188 37176 8192
rect 37112 8132 37116 8188
rect 37116 8132 37172 8188
rect 37172 8132 37176 8188
rect 37112 8128 37176 8132
rect 37192 8188 37256 8192
rect 37192 8132 37196 8188
rect 37196 8132 37252 8188
rect 37252 8132 37256 8188
rect 37192 8128 37256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 7612 7644 7676 7648
rect 7612 7588 7616 7644
rect 7616 7588 7672 7644
rect 7672 7588 7676 7644
rect 7612 7584 7676 7588
rect 7692 7644 7756 7648
rect 7692 7588 7696 7644
rect 7696 7588 7752 7644
rect 7752 7588 7756 7644
rect 7692 7584 7756 7588
rect 7772 7644 7836 7648
rect 7772 7588 7776 7644
rect 7776 7588 7832 7644
rect 7832 7588 7836 7644
rect 7772 7584 7836 7588
rect 7852 7644 7916 7648
rect 7852 7588 7856 7644
rect 7856 7588 7912 7644
rect 7912 7588 7916 7644
rect 7852 7584 7916 7588
rect 12612 7644 12676 7648
rect 12612 7588 12616 7644
rect 12616 7588 12672 7644
rect 12672 7588 12676 7644
rect 12612 7584 12676 7588
rect 12692 7644 12756 7648
rect 12692 7588 12696 7644
rect 12696 7588 12752 7644
rect 12752 7588 12756 7644
rect 12692 7584 12756 7588
rect 12772 7644 12836 7648
rect 12772 7588 12776 7644
rect 12776 7588 12832 7644
rect 12832 7588 12836 7644
rect 12772 7584 12836 7588
rect 12852 7644 12916 7648
rect 12852 7588 12856 7644
rect 12856 7588 12912 7644
rect 12912 7588 12916 7644
rect 12852 7584 12916 7588
rect 17612 7644 17676 7648
rect 17612 7588 17616 7644
rect 17616 7588 17672 7644
rect 17672 7588 17676 7644
rect 17612 7584 17676 7588
rect 17692 7644 17756 7648
rect 17692 7588 17696 7644
rect 17696 7588 17752 7644
rect 17752 7588 17756 7644
rect 17692 7584 17756 7588
rect 17772 7644 17836 7648
rect 17772 7588 17776 7644
rect 17776 7588 17832 7644
rect 17832 7588 17836 7644
rect 17772 7584 17836 7588
rect 17852 7644 17916 7648
rect 17852 7588 17856 7644
rect 17856 7588 17912 7644
rect 17912 7588 17916 7644
rect 17852 7584 17916 7588
rect 22612 7644 22676 7648
rect 22612 7588 22616 7644
rect 22616 7588 22672 7644
rect 22672 7588 22676 7644
rect 22612 7584 22676 7588
rect 22692 7644 22756 7648
rect 22692 7588 22696 7644
rect 22696 7588 22752 7644
rect 22752 7588 22756 7644
rect 22692 7584 22756 7588
rect 22772 7644 22836 7648
rect 22772 7588 22776 7644
rect 22776 7588 22832 7644
rect 22832 7588 22836 7644
rect 22772 7584 22836 7588
rect 22852 7644 22916 7648
rect 22852 7588 22856 7644
rect 22856 7588 22912 7644
rect 22912 7588 22916 7644
rect 22852 7584 22916 7588
rect 27612 7644 27676 7648
rect 27612 7588 27616 7644
rect 27616 7588 27672 7644
rect 27672 7588 27676 7644
rect 27612 7584 27676 7588
rect 27692 7644 27756 7648
rect 27692 7588 27696 7644
rect 27696 7588 27752 7644
rect 27752 7588 27756 7644
rect 27692 7584 27756 7588
rect 27772 7644 27836 7648
rect 27772 7588 27776 7644
rect 27776 7588 27832 7644
rect 27832 7588 27836 7644
rect 27772 7584 27836 7588
rect 27852 7644 27916 7648
rect 27852 7588 27856 7644
rect 27856 7588 27912 7644
rect 27912 7588 27916 7644
rect 27852 7584 27916 7588
rect 32612 7644 32676 7648
rect 32612 7588 32616 7644
rect 32616 7588 32672 7644
rect 32672 7588 32676 7644
rect 32612 7584 32676 7588
rect 32692 7644 32756 7648
rect 32692 7588 32696 7644
rect 32696 7588 32752 7644
rect 32752 7588 32756 7644
rect 32692 7584 32756 7588
rect 32772 7644 32836 7648
rect 32772 7588 32776 7644
rect 32776 7588 32832 7644
rect 32832 7588 32836 7644
rect 32772 7584 32836 7588
rect 32852 7644 32916 7648
rect 32852 7588 32856 7644
rect 32856 7588 32912 7644
rect 32912 7588 32916 7644
rect 32852 7584 32916 7588
rect 37612 7644 37676 7648
rect 37612 7588 37616 7644
rect 37616 7588 37672 7644
rect 37672 7588 37676 7644
rect 37612 7584 37676 7588
rect 37692 7644 37756 7648
rect 37692 7588 37696 7644
rect 37696 7588 37752 7644
rect 37752 7588 37756 7644
rect 37692 7584 37756 7588
rect 37772 7644 37836 7648
rect 37772 7588 37776 7644
rect 37776 7588 37832 7644
rect 37832 7588 37836 7644
rect 37772 7584 37836 7588
rect 37852 7644 37916 7648
rect 37852 7588 37856 7644
rect 37856 7588 37912 7644
rect 37912 7588 37916 7644
rect 37852 7584 37916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 6952 7100 7016 7104
rect 6952 7044 6956 7100
rect 6956 7044 7012 7100
rect 7012 7044 7016 7100
rect 6952 7040 7016 7044
rect 7032 7100 7096 7104
rect 7032 7044 7036 7100
rect 7036 7044 7092 7100
rect 7092 7044 7096 7100
rect 7032 7040 7096 7044
rect 7112 7100 7176 7104
rect 7112 7044 7116 7100
rect 7116 7044 7172 7100
rect 7172 7044 7176 7100
rect 7112 7040 7176 7044
rect 7192 7100 7256 7104
rect 7192 7044 7196 7100
rect 7196 7044 7252 7100
rect 7252 7044 7256 7100
rect 7192 7040 7256 7044
rect 11952 7100 12016 7104
rect 11952 7044 11956 7100
rect 11956 7044 12012 7100
rect 12012 7044 12016 7100
rect 11952 7040 12016 7044
rect 12032 7100 12096 7104
rect 12032 7044 12036 7100
rect 12036 7044 12092 7100
rect 12092 7044 12096 7100
rect 12032 7040 12096 7044
rect 12112 7100 12176 7104
rect 12112 7044 12116 7100
rect 12116 7044 12172 7100
rect 12172 7044 12176 7100
rect 12112 7040 12176 7044
rect 12192 7100 12256 7104
rect 12192 7044 12196 7100
rect 12196 7044 12252 7100
rect 12252 7044 12256 7100
rect 12192 7040 12256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 21952 7100 22016 7104
rect 21952 7044 21956 7100
rect 21956 7044 22012 7100
rect 22012 7044 22016 7100
rect 21952 7040 22016 7044
rect 22032 7100 22096 7104
rect 22032 7044 22036 7100
rect 22036 7044 22092 7100
rect 22092 7044 22096 7100
rect 22032 7040 22096 7044
rect 22112 7100 22176 7104
rect 22112 7044 22116 7100
rect 22116 7044 22172 7100
rect 22172 7044 22176 7100
rect 22112 7040 22176 7044
rect 22192 7100 22256 7104
rect 22192 7044 22196 7100
rect 22196 7044 22252 7100
rect 22252 7044 22256 7100
rect 22192 7040 22256 7044
rect 26952 7100 27016 7104
rect 26952 7044 26956 7100
rect 26956 7044 27012 7100
rect 27012 7044 27016 7100
rect 26952 7040 27016 7044
rect 27032 7100 27096 7104
rect 27032 7044 27036 7100
rect 27036 7044 27092 7100
rect 27092 7044 27096 7100
rect 27032 7040 27096 7044
rect 27112 7100 27176 7104
rect 27112 7044 27116 7100
rect 27116 7044 27172 7100
rect 27172 7044 27176 7100
rect 27112 7040 27176 7044
rect 27192 7100 27256 7104
rect 27192 7044 27196 7100
rect 27196 7044 27252 7100
rect 27252 7044 27256 7100
rect 27192 7040 27256 7044
rect 31952 7100 32016 7104
rect 31952 7044 31956 7100
rect 31956 7044 32012 7100
rect 32012 7044 32016 7100
rect 31952 7040 32016 7044
rect 32032 7100 32096 7104
rect 32032 7044 32036 7100
rect 32036 7044 32092 7100
rect 32092 7044 32096 7100
rect 32032 7040 32096 7044
rect 32112 7100 32176 7104
rect 32112 7044 32116 7100
rect 32116 7044 32172 7100
rect 32172 7044 32176 7100
rect 32112 7040 32176 7044
rect 32192 7100 32256 7104
rect 32192 7044 32196 7100
rect 32196 7044 32252 7100
rect 32252 7044 32256 7100
rect 32192 7040 32256 7044
rect 36952 7100 37016 7104
rect 36952 7044 36956 7100
rect 36956 7044 37012 7100
rect 37012 7044 37016 7100
rect 36952 7040 37016 7044
rect 37032 7100 37096 7104
rect 37032 7044 37036 7100
rect 37036 7044 37092 7100
rect 37092 7044 37096 7100
rect 37032 7040 37096 7044
rect 37112 7100 37176 7104
rect 37112 7044 37116 7100
rect 37116 7044 37172 7100
rect 37172 7044 37176 7100
rect 37112 7040 37176 7044
rect 37192 7100 37256 7104
rect 37192 7044 37196 7100
rect 37196 7044 37252 7100
rect 37252 7044 37256 7100
rect 37192 7040 37256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 7612 6556 7676 6560
rect 7612 6500 7616 6556
rect 7616 6500 7672 6556
rect 7672 6500 7676 6556
rect 7612 6496 7676 6500
rect 7692 6556 7756 6560
rect 7692 6500 7696 6556
rect 7696 6500 7752 6556
rect 7752 6500 7756 6556
rect 7692 6496 7756 6500
rect 7772 6556 7836 6560
rect 7772 6500 7776 6556
rect 7776 6500 7832 6556
rect 7832 6500 7836 6556
rect 7772 6496 7836 6500
rect 7852 6556 7916 6560
rect 7852 6500 7856 6556
rect 7856 6500 7912 6556
rect 7912 6500 7916 6556
rect 7852 6496 7916 6500
rect 12612 6556 12676 6560
rect 12612 6500 12616 6556
rect 12616 6500 12672 6556
rect 12672 6500 12676 6556
rect 12612 6496 12676 6500
rect 12692 6556 12756 6560
rect 12692 6500 12696 6556
rect 12696 6500 12752 6556
rect 12752 6500 12756 6556
rect 12692 6496 12756 6500
rect 12772 6556 12836 6560
rect 12772 6500 12776 6556
rect 12776 6500 12832 6556
rect 12832 6500 12836 6556
rect 12772 6496 12836 6500
rect 12852 6556 12916 6560
rect 12852 6500 12856 6556
rect 12856 6500 12912 6556
rect 12912 6500 12916 6556
rect 12852 6496 12916 6500
rect 17612 6556 17676 6560
rect 17612 6500 17616 6556
rect 17616 6500 17672 6556
rect 17672 6500 17676 6556
rect 17612 6496 17676 6500
rect 17692 6556 17756 6560
rect 17692 6500 17696 6556
rect 17696 6500 17752 6556
rect 17752 6500 17756 6556
rect 17692 6496 17756 6500
rect 17772 6556 17836 6560
rect 17772 6500 17776 6556
rect 17776 6500 17832 6556
rect 17832 6500 17836 6556
rect 17772 6496 17836 6500
rect 17852 6556 17916 6560
rect 17852 6500 17856 6556
rect 17856 6500 17912 6556
rect 17912 6500 17916 6556
rect 17852 6496 17916 6500
rect 22612 6556 22676 6560
rect 22612 6500 22616 6556
rect 22616 6500 22672 6556
rect 22672 6500 22676 6556
rect 22612 6496 22676 6500
rect 22692 6556 22756 6560
rect 22692 6500 22696 6556
rect 22696 6500 22752 6556
rect 22752 6500 22756 6556
rect 22692 6496 22756 6500
rect 22772 6556 22836 6560
rect 22772 6500 22776 6556
rect 22776 6500 22832 6556
rect 22832 6500 22836 6556
rect 22772 6496 22836 6500
rect 22852 6556 22916 6560
rect 22852 6500 22856 6556
rect 22856 6500 22912 6556
rect 22912 6500 22916 6556
rect 22852 6496 22916 6500
rect 27612 6556 27676 6560
rect 27612 6500 27616 6556
rect 27616 6500 27672 6556
rect 27672 6500 27676 6556
rect 27612 6496 27676 6500
rect 27692 6556 27756 6560
rect 27692 6500 27696 6556
rect 27696 6500 27752 6556
rect 27752 6500 27756 6556
rect 27692 6496 27756 6500
rect 27772 6556 27836 6560
rect 27772 6500 27776 6556
rect 27776 6500 27832 6556
rect 27832 6500 27836 6556
rect 27772 6496 27836 6500
rect 27852 6556 27916 6560
rect 27852 6500 27856 6556
rect 27856 6500 27912 6556
rect 27912 6500 27916 6556
rect 27852 6496 27916 6500
rect 32612 6556 32676 6560
rect 32612 6500 32616 6556
rect 32616 6500 32672 6556
rect 32672 6500 32676 6556
rect 32612 6496 32676 6500
rect 32692 6556 32756 6560
rect 32692 6500 32696 6556
rect 32696 6500 32752 6556
rect 32752 6500 32756 6556
rect 32692 6496 32756 6500
rect 32772 6556 32836 6560
rect 32772 6500 32776 6556
rect 32776 6500 32832 6556
rect 32832 6500 32836 6556
rect 32772 6496 32836 6500
rect 32852 6556 32916 6560
rect 32852 6500 32856 6556
rect 32856 6500 32912 6556
rect 32912 6500 32916 6556
rect 32852 6496 32916 6500
rect 37612 6556 37676 6560
rect 37612 6500 37616 6556
rect 37616 6500 37672 6556
rect 37672 6500 37676 6556
rect 37612 6496 37676 6500
rect 37692 6556 37756 6560
rect 37692 6500 37696 6556
rect 37696 6500 37752 6556
rect 37752 6500 37756 6556
rect 37692 6496 37756 6500
rect 37772 6556 37836 6560
rect 37772 6500 37776 6556
rect 37776 6500 37832 6556
rect 37832 6500 37836 6556
rect 37772 6496 37836 6500
rect 37852 6556 37916 6560
rect 37852 6500 37856 6556
rect 37856 6500 37912 6556
rect 37912 6500 37916 6556
rect 37852 6496 37916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 6952 6012 7016 6016
rect 6952 5956 6956 6012
rect 6956 5956 7012 6012
rect 7012 5956 7016 6012
rect 6952 5952 7016 5956
rect 7032 6012 7096 6016
rect 7032 5956 7036 6012
rect 7036 5956 7092 6012
rect 7092 5956 7096 6012
rect 7032 5952 7096 5956
rect 7112 6012 7176 6016
rect 7112 5956 7116 6012
rect 7116 5956 7172 6012
rect 7172 5956 7176 6012
rect 7112 5952 7176 5956
rect 7192 6012 7256 6016
rect 7192 5956 7196 6012
rect 7196 5956 7252 6012
rect 7252 5956 7256 6012
rect 7192 5952 7256 5956
rect 11952 6012 12016 6016
rect 11952 5956 11956 6012
rect 11956 5956 12012 6012
rect 12012 5956 12016 6012
rect 11952 5952 12016 5956
rect 12032 6012 12096 6016
rect 12032 5956 12036 6012
rect 12036 5956 12092 6012
rect 12092 5956 12096 6012
rect 12032 5952 12096 5956
rect 12112 6012 12176 6016
rect 12112 5956 12116 6012
rect 12116 5956 12172 6012
rect 12172 5956 12176 6012
rect 12112 5952 12176 5956
rect 12192 6012 12256 6016
rect 12192 5956 12196 6012
rect 12196 5956 12252 6012
rect 12252 5956 12256 6012
rect 12192 5952 12256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 21952 6012 22016 6016
rect 21952 5956 21956 6012
rect 21956 5956 22012 6012
rect 22012 5956 22016 6012
rect 21952 5952 22016 5956
rect 22032 6012 22096 6016
rect 22032 5956 22036 6012
rect 22036 5956 22092 6012
rect 22092 5956 22096 6012
rect 22032 5952 22096 5956
rect 22112 6012 22176 6016
rect 22112 5956 22116 6012
rect 22116 5956 22172 6012
rect 22172 5956 22176 6012
rect 22112 5952 22176 5956
rect 22192 6012 22256 6016
rect 22192 5956 22196 6012
rect 22196 5956 22252 6012
rect 22252 5956 22256 6012
rect 22192 5952 22256 5956
rect 26952 6012 27016 6016
rect 26952 5956 26956 6012
rect 26956 5956 27012 6012
rect 27012 5956 27016 6012
rect 26952 5952 27016 5956
rect 27032 6012 27096 6016
rect 27032 5956 27036 6012
rect 27036 5956 27092 6012
rect 27092 5956 27096 6012
rect 27032 5952 27096 5956
rect 27112 6012 27176 6016
rect 27112 5956 27116 6012
rect 27116 5956 27172 6012
rect 27172 5956 27176 6012
rect 27112 5952 27176 5956
rect 27192 6012 27256 6016
rect 27192 5956 27196 6012
rect 27196 5956 27252 6012
rect 27252 5956 27256 6012
rect 27192 5952 27256 5956
rect 31952 6012 32016 6016
rect 31952 5956 31956 6012
rect 31956 5956 32012 6012
rect 32012 5956 32016 6012
rect 31952 5952 32016 5956
rect 32032 6012 32096 6016
rect 32032 5956 32036 6012
rect 32036 5956 32092 6012
rect 32092 5956 32096 6012
rect 32032 5952 32096 5956
rect 32112 6012 32176 6016
rect 32112 5956 32116 6012
rect 32116 5956 32172 6012
rect 32172 5956 32176 6012
rect 32112 5952 32176 5956
rect 32192 6012 32256 6016
rect 32192 5956 32196 6012
rect 32196 5956 32252 6012
rect 32252 5956 32256 6012
rect 32192 5952 32256 5956
rect 36952 6012 37016 6016
rect 36952 5956 36956 6012
rect 36956 5956 37012 6012
rect 37012 5956 37016 6012
rect 36952 5952 37016 5956
rect 37032 6012 37096 6016
rect 37032 5956 37036 6012
rect 37036 5956 37092 6012
rect 37092 5956 37096 6012
rect 37032 5952 37096 5956
rect 37112 6012 37176 6016
rect 37112 5956 37116 6012
rect 37116 5956 37172 6012
rect 37172 5956 37176 6012
rect 37112 5952 37176 5956
rect 37192 6012 37256 6016
rect 37192 5956 37196 6012
rect 37196 5956 37252 6012
rect 37252 5956 37256 6012
rect 37192 5952 37256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 7612 5468 7676 5472
rect 7612 5412 7616 5468
rect 7616 5412 7672 5468
rect 7672 5412 7676 5468
rect 7612 5408 7676 5412
rect 7692 5468 7756 5472
rect 7692 5412 7696 5468
rect 7696 5412 7752 5468
rect 7752 5412 7756 5468
rect 7692 5408 7756 5412
rect 7772 5468 7836 5472
rect 7772 5412 7776 5468
rect 7776 5412 7832 5468
rect 7832 5412 7836 5468
rect 7772 5408 7836 5412
rect 7852 5468 7916 5472
rect 7852 5412 7856 5468
rect 7856 5412 7912 5468
rect 7912 5412 7916 5468
rect 7852 5408 7916 5412
rect 12612 5468 12676 5472
rect 12612 5412 12616 5468
rect 12616 5412 12672 5468
rect 12672 5412 12676 5468
rect 12612 5408 12676 5412
rect 12692 5468 12756 5472
rect 12692 5412 12696 5468
rect 12696 5412 12752 5468
rect 12752 5412 12756 5468
rect 12692 5408 12756 5412
rect 12772 5468 12836 5472
rect 12772 5412 12776 5468
rect 12776 5412 12832 5468
rect 12832 5412 12836 5468
rect 12772 5408 12836 5412
rect 12852 5468 12916 5472
rect 12852 5412 12856 5468
rect 12856 5412 12912 5468
rect 12912 5412 12916 5468
rect 12852 5408 12916 5412
rect 17612 5468 17676 5472
rect 17612 5412 17616 5468
rect 17616 5412 17672 5468
rect 17672 5412 17676 5468
rect 17612 5408 17676 5412
rect 17692 5468 17756 5472
rect 17692 5412 17696 5468
rect 17696 5412 17752 5468
rect 17752 5412 17756 5468
rect 17692 5408 17756 5412
rect 17772 5468 17836 5472
rect 17772 5412 17776 5468
rect 17776 5412 17832 5468
rect 17832 5412 17836 5468
rect 17772 5408 17836 5412
rect 17852 5468 17916 5472
rect 17852 5412 17856 5468
rect 17856 5412 17912 5468
rect 17912 5412 17916 5468
rect 17852 5408 17916 5412
rect 22612 5468 22676 5472
rect 22612 5412 22616 5468
rect 22616 5412 22672 5468
rect 22672 5412 22676 5468
rect 22612 5408 22676 5412
rect 22692 5468 22756 5472
rect 22692 5412 22696 5468
rect 22696 5412 22752 5468
rect 22752 5412 22756 5468
rect 22692 5408 22756 5412
rect 22772 5468 22836 5472
rect 22772 5412 22776 5468
rect 22776 5412 22832 5468
rect 22832 5412 22836 5468
rect 22772 5408 22836 5412
rect 22852 5468 22916 5472
rect 22852 5412 22856 5468
rect 22856 5412 22912 5468
rect 22912 5412 22916 5468
rect 22852 5408 22916 5412
rect 27612 5468 27676 5472
rect 27612 5412 27616 5468
rect 27616 5412 27672 5468
rect 27672 5412 27676 5468
rect 27612 5408 27676 5412
rect 27692 5468 27756 5472
rect 27692 5412 27696 5468
rect 27696 5412 27752 5468
rect 27752 5412 27756 5468
rect 27692 5408 27756 5412
rect 27772 5468 27836 5472
rect 27772 5412 27776 5468
rect 27776 5412 27832 5468
rect 27832 5412 27836 5468
rect 27772 5408 27836 5412
rect 27852 5468 27916 5472
rect 27852 5412 27856 5468
rect 27856 5412 27912 5468
rect 27912 5412 27916 5468
rect 27852 5408 27916 5412
rect 32612 5468 32676 5472
rect 32612 5412 32616 5468
rect 32616 5412 32672 5468
rect 32672 5412 32676 5468
rect 32612 5408 32676 5412
rect 32692 5468 32756 5472
rect 32692 5412 32696 5468
rect 32696 5412 32752 5468
rect 32752 5412 32756 5468
rect 32692 5408 32756 5412
rect 32772 5468 32836 5472
rect 32772 5412 32776 5468
rect 32776 5412 32832 5468
rect 32832 5412 32836 5468
rect 32772 5408 32836 5412
rect 32852 5468 32916 5472
rect 32852 5412 32856 5468
rect 32856 5412 32912 5468
rect 32912 5412 32916 5468
rect 32852 5408 32916 5412
rect 37612 5468 37676 5472
rect 37612 5412 37616 5468
rect 37616 5412 37672 5468
rect 37672 5412 37676 5468
rect 37612 5408 37676 5412
rect 37692 5468 37756 5472
rect 37692 5412 37696 5468
rect 37696 5412 37752 5468
rect 37752 5412 37756 5468
rect 37692 5408 37756 5412
rect 37772 5468 37836 5472
rect 37772 5412 37776 5468
rect 37776 5412 37832 5468
rect 37832 5412 37836 5468
rect 37772 5408 37836 5412
rect 37852 5468 37916 5472
rect 37852 5412 37856 5468
rect 37856 5412 37912 5468
rect 37912 5412 37916 5468
rect 37852 5408 37916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 6952 4924 7016 4928
rect 6952 4868 6956 4924
rect 6956 4868 7012 4924
rect 7012 4868 7016 4924
rect 6952 4864 7016 4868
rect 7032 4924 7096 4928
rect 7032 4868 7036 4924
rect 7036 4868 7092 4924
rect 7092 4868 7096 4924
rect 7032 4864 7096 4868
rect 7112 4924 7176 4928
rect 7112 4868 7116 4924
rect 7116 4868 7172 4924
rect 7172 4868 7176 4924
rect 7112 4864 7176 4868
rect 7192 4924 7256 4928
rect 7192 4868 7196 4924
rect 7196 4868 7252 4924
rect 7252 4868 7256 4924
rect 7192 4864 7256 4868
rect 11952 4924 12016 4928
rect 11952 4868 11956 4924
rect 11956 4868 12012 4924
rect 12012 4868 12016 4924
rect 11952 4864 12016 4868
rect 12032 4924 12096 4928
rect 12032 4868 12036 4924
rect 12036 4868 12092 4924
rect 12092 4868 12096 4924
rect 12032 4864 12096 4868
rect 12112 4924 12176 4928
rect 12112 4868 12116 4924
rect 12116 4868 12172 4924
rect 12172 4868 12176 4924
rect 12112 4864 12176 4868
rect 12192 4924 12256 4928
rect 12192 4868 12196 4924
rect 12196 4868 12252 4924
rect 12252 4868 12256 4924
rect 12192 4864 12256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 21952 4924 22016 4928
rect 21952 4868 21956 4924
rect 21956 4868 22012 4924
rect 22012 4868 22016 4924
rect 21952 4864 22016 4868
rect 22032 4924 22096 4928
rect 22032 4868 22036 4924
rect 22036 4868 22092 4924
rect 22092 4868 22096 4924
rect 22032 4864 22096 4868
rect 22112 4924 22176 4928
rect 22112 4868 22116 4924
rect 22116 4868 22172 4924
rect 22172 4868 22176 4924
rect 22112 4864 22176 4868
rect 22192 4924 22256 4928
rect 22192 4868 22196 4924
rect 22196 4868 22252 4924
rect 22252 4868 22256 4924
rect 22192 4864 22256 4868
rect 26952 4924 27016 4928
rect 26952 4868 26956 4924
rect 26956 4868 27012 4924
rect 27012 4868 27016 4924
rect 26952 4864 27016 4868
rect 27032 4924 27096 4928
rect 27032 4868 27036 4924
rect 27036 4868 27092 4924
rect 27092 4868 27096 4924
rect 27032 4864 27096 4868
rect 27112 4924 27176 4928
rect 27112 4868 27116 4924
rect 27116 4868 27172 4924
rect 27172 4868 27176 4924
rect 27112 4864 27176 4868
rect 27192 4924 27256 4928
rect 27192 4868 27196 4924
rect 27196 4868 27252 4924
rect 27252 4868 27256 4924
rect 27192 4864 27256 4868
rect 31952 4924 32016 4928
rect 31952 4868 31956 4924
rect 31956 4868 32012 4924
rect 32012 4868 32016 4924
rect 31952 4864 32016 4868
rect 32032 4924 32096 4928
rect 32032 4868 32036 4924
rect 32036 4868 32092 4924
rect 32092 4868 32096 4924
rect 32032 4864 32096 4868
rect 32112 4924 32176 4928
rect 32112 4868 32116 4924
rect 32116 4868 32172 4924
rect 32172 4868 32176 4924
rect 32112 4864 32176 4868
rect 32192 4924 32256 4928
rect 32192 4868 32196 4924
rect 32196 4868 32252 4924
rect 32252 4868 32256 4924
rect 32192 4864 32256 4868
rect 36952 4924 37016 4928
rect 36952 4868 36956 4924
rect 36956 4868 37012 4924
rect 37012 4868 37016 4924
rect 36952 4864 37016 4868
rect 37032 4924 37096 4928
rect 37032 4868 37036 4924
rect 37036 4868 37092 4924
rect 37092 4868 37096 4924
rect 37032 4864 37096 4868
rect 37112 4924 37176 4928
rect 37112 4868 37116 4924
rect 37116 4868 37172 4924
rect 37172 4868 37176 4924
rect 37112 4864 37176 4868
rect 37192 4924 37256 4928
rect 37192 4868 37196 4924
rect 37196 4868 37252 4924
rect 37252 4868 37256 4924
rect 37192 4864 37256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 7612 4380 7676 4384
rect 7612 4324 7616 4380
rect 7616 4324 7672 4380
rect 7672 4324 7676 4380
rect 7612 4320 7676 4324
rect 7692 4380 7756 4384
rect 7692 4324 7696 4380
rect 7696 4324 7752 4380
rect 7752 4324 7756 4380
rect 7692 4320 7756 4324
rect 7772 4380 7836 4384
rect 7772 4324 7776 4380
rect 7776 4324 7832 4380
rect 7832 4324 7836 4380
rect 7772 4320 7836 4324
rect 7852 4380 7916 4384
rect 7852 4324 7856 4380
rect 7856 4324 7912 4380
rect 7912 4324 7916 4380
rect 7852 4320 7916 4324
rect 12612 4380 12676 4384
rect 12612 4324 12616 4380
rect 12616 4324 12672 4380
rect 12672 4324 12676 4380
rect 12612 4320 12676 4324
rect 12692 4380 12756 4384
rect 12692 4324 12696 4380
rect 12696 4324 12752 4380
rect 12752 4324 12756 4380
rect 12692 4320 12756 4324
rect 12772 4380 12836 4384
rect 12772 4324 12776 4380
rect 12776 4324 12832 4380
rect 12832 4324 12836 4380
rect 12772 4320 12836 4324
rect 12852 4380 12916 4384
rect 12852 4324 12856 4380
rect 12856 4324 12912 4380
rect 12912 4324 12916 4380
rect 12852 4320 12916 4324
rect 17612 4380 17676 4384
rect 17612 4324 17616 4380
rect 17616 4324 17672 4380
rect 17672 4324 17676 4380
rect 17612 4320 17676 4324
rect 17692 4380 17756 4384
rect 17692 4324 17696 4380
rect 17696 4324 17752 4380
rect 17752 4324 17756 4380
rect 17692 4320 17756 4324
rect 17772 4380 17836 4384
rect 17772 4324 17776 4380
rect 17776 4324 17832 4380
rect 17832 4324 17836 4380
rect 17772 4320 17836 4324
rect 17852 4380 17916 4384
rect 17852 4324 17856 4380
rect 17856 4324 17912 4380
rect 17912 4324 17916 4380
rect 17852 4320 17916 4324
rect 22612 4380 22676 4384
rect 22612 4324 22616 4380
rect 22616 4324 22672 4380
rect 22672 4324 22676 4380
rect 22612 4320 22676 4324
rect 22692 4380 22756 4384
rect 22692 4324 22696 4380
rect 22696 4324 22752 4380
rect 22752 4324 22756 4380
rect 22692 4320 22756 4324
rect 22772 4380 22836 4384
rect 22772 4324 22776 4380
rect 22776 4324 22832 4380
rect 22832 4324 22836 4380
rect 22772 4320 22836 4324
rect 22852 4380 22916 4384
rect 22852 4324 22856 4380
rect 22856 4324 22912 4380
rect 22912 4324 22916 4380
rect 22852 4320 22916 4324
rect 27612 4380 27676 4384
rect 27612 4324 27616 4380
rect 27616 4324 27672 4380
rect 27672 4324 27676 4380
rect 27612 4320 27676 4324
rect 27692 4380 27756 4384
rect 27692 4324 27696 4380
rect 27696 4324 27752 4380
rect 27752 4324 27756 4380
rect 27692 4320 27756 4324
rect 27772 4380 27836 4384
rect 27772 4324 27776 4380
rect 27776 4324 27832 4380
rect 27832 4324 27836 4380
rect 27772 4320 27836 4324
rect 27852 4380 27916 4384
rect 27852 4324 27856 4380
rect 27856 4324 27912 4380
rect 27912 4324 27916 4380
rect 27852 4320 27916 4324
rect 32612 4380 32676 4384
rect 32612 4324 32616 4380
rect 32616 4324 32672 4380
rect 32672 4324 32676 4380
rect 32612 4320 32676 4324
rect 32692 4380 32756 4384
rect 32692 4324 32696 4380
rect 32696 4324 32752 4380
rect 32752 4324 32756 4380
rect 32692 4320 32756 4324
rect 32772 4380 32836 4384
rect 32772 4324 32776 4380
rect 32776 4324 32832 4380
rect 32832 4324 32836 4380
rect 32772 4320 32836 4324
rect 32852 4380 32916 4384
rect 32852 4324 32856 4380
rect 32856 4324 32912 4380
rect 32912 4324 32916 4380
rect 32852 4320 32916 4324
rect 37612 4380 37676 4384
rect 37612 4324 37616 4380
rect 37616 4324 37672 4380
rect 37672 4324 37676 4380
rect 37612 4320 37676 4324
rect 37692 4380 37756 4384
rect 37692 4324 37696 4380
rect 37696 4324 37752 4380
rect 37752 4324 37756 4380
rect 37692 4320 37756 4324
rect 37772 4380 37836 4384
rect 37772 4324 37776 4380
rect 37776 4324 37832 4380
rect 37832 4324 37836 4380
rect 37772 4320 37836 4324
rect 37852 4380 37916 4384
rect 37852 4324 37856 4380
rect 37856 4324 37912 4380
rect 37912 4324 37916 4380
rect 37852 4320 37916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 6952 3836 7016 3840
rect 6952 3780 6956 3836
rect 6956 3780 7012 3836
rect 7012 3780 7016 3836
rect 6952 3776 7016 3780
rect 7032 3836 7096 3840
rect 7032 3780 7036 3836
rect 7036 3780 7092 3836
rect 7092 3780 7096 3836
rect 7032 3776 7096 3780
rect 7112 3836 7176 3840
rect 7112 3780 7116 3836
rect 7116 3780 7172 3836
rect 7172 3780 7176 3836
rect 7112 3776 7176 3780
rect 7192 3836 7256 3840
rect 7192 3780 7196 3836
rect 7196 3780 7252 3836
rect 7252 3780 7256 3836
rect 7192 3776 7256 3780
rect 11952 3836 12016 3840
rect 11952 3780 11956 3836
rect 11956 3780 12012 3836
rect 12012 3780 12016 3836
rect 11952 3776 12016 3780
rect 12032 3836 12096 3840
rect 12032 3780 12036 3836
rect 12036 3780 12092 3836
rect 12092 3780 12096 3836
rect 12032 3776 12096 3780
rect 12112 3836 12176 3840
rect 12112 3780 12116 3836
rect 12116 3780 12172 3836
rect 12172 3780 12176 3836
rect 12112 3776 12176 3780
rect 12192 3836 12256 3840
rect 12192 3780 12196 3836
rect 12196 3780 12252 3836
rect 12252 3780 12256 3836
rect 12192 3776 12256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 21952 3836 22016 3840
rect 21952 3780 21956 3836
rect 21956 3780 22012 3836
rect 22012 3780 22016 3836
rect 21952 3776 22016 3780
rect 22032 3836 22096 3840
rect 22032 3780 22036 3836
rect 22036 3780 22092 3836
rect 22092 3780 22096 3836
rect 22032 3776 22096 3780
rect 22112 3836 22176 3840
rect 22112 3780 22116 3836
rect 22116 3780 22172 3836
rect 22172 3780 22176 3836
rect 22112 3776 22176 3780
rect 22192 3836 22256 3840
rect 22192 3780 22196 3836
rect 22196 3780 22252 3836
rect 22252 3780 22256 3836
rect 22192 3776 22256 3780
rect 26952 3836 27016 3840
rect 26952 3780 26956 3836
rect 26956 3780 27012 3836
rect 27012 3780 27016 3836
rect 26952 3776 27016 3780
rect 27032 3836 27096 3840
rect 27032 3780 27036 3836
rect 27036 3780 27092 3836
rect 27092 3780 27096 3836
rect 27032 3776 27096 3780
rect 27112 3836 27176 3840
rect 27112 3780 27116 3836
rect 27116 3780 27172 3836
rect 27172 3780 27176 3836
rect 27112 3776 27176 3780
rect 27192 3836 27256 3840
rect 27192 3780 27196 3836
rect 27196 3780 27252 3836
rect 27252 3780 27256 3836
rect 27192 3776 27256 3780
rect 31952 3836 32016 3840
rect 31952 3780 31956 3836
rect 31956 3780 32012 3836
rect 32012 3780 32016 3836
rect 31952 3776 32016 3780
rect 32032 3836 32096 3840
rect 32032 3780 32036 3836
rect 32036 3780 32092 3836
rect 32092 3780 32096 3836
rect 32032 3776 32096 3780
rect 32112 3836 32176 3840
rect 32112 3780 32116 3836
rect 32116 3780 32172 3836
rect 32172 3780 32176 3836
rect 32112 3776 32176 3780
rect 32192 3836 32256 3840
rect 32192 3780 32196 3836
rect 32196 3780 32252 3836
rect 32252 3780 32256 3836
rect 32192 3776 32256 3780
rect 36952 3836 37016 3840
rect 36952 3780 36956 3836
rect 36956 3780 37012 3836
rect 37012 3780 37016 3836
rect 36952 3776 37016 3780
rect 37032 3836 37096 3840
rect 37032 3780 37036 3836
rect 37036 3780 37092 3836
rect 37092 3780 37096 3836
rect 37032 3776 37096 3780
rect 37112 3836 37176 3840
rect 37112 3780 37116 3836
rect 37116 3780 37172 3836
rect 37172 3780 37176 3836
rect 37112 3776 37176 3780
rect 37192 3836 37256 3840
rect 37192 3780 37196 3836
rect 37196 3780 37252 3836
rect 37252 3780 37256 3836
rect 37192 3776 37256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 7612 3292 7676 3296
rect 7612 3236 7616 3292
rect 7616 3236 7672 3292
rect 7672 3236 7676 3292
rect 7612 3232 7676 3236
rect 7692 3292 7756 3296
rect 7692 3236 7696 3292
rect 7696 3236 7752 3292
rect 7752 3236 7756 3292
rect 7692 3232 7756 3236
rect 7772 3292 7836 3296
rect 7772 3236 7776 3292
rect 7776 3236 7832 3292
rect 7832 3236 7836 3292
rect 7772 3232 7836 3236
rect 7852 3292 7916 3296
rect 7852 3236 7856 3292
rect 7856 3236 7912 3292
rect 7912 3236 7916 3292
rect 7852 3232 7916 3236
rect 12612 3292 12676 3296
rect 12612 3236 12616 3292
rect 12616 3236 12672 3292
rect 12672 3236 12676 3292
rect 12612 3232 12676 3236
rect 12692 3292 12756 3296
rect 12692 3236 12696 3292
rect 12696 3236 12752 3292
rect 12752 3236 12756 3292
rect 12692 3232 12756 3236
rect 12772 3292 12836 3296
rect 12772 3236 12776 3292
rect 12776 3236 12832 3292
rect 12832 3236 12836 3292
rect 12772 3232 12836 3236
rect 12852 3292 12916 3296
rect 12852 3236 12856 3292
rect 12856 3236 12912 3292
rect 12912 3236 12916 3292
rect 12852 3232 12916 3236
rect 17612 3292 17676 3296
rect 17612 3236 17616 3292
rect 17616 3236 17672 3292
rect 17672 3236 17676 3292
rect 17612 3232 17676 3236
rect 17692 3292 17756 3296
rect 17692 3236 17696 3292
rect 17696 3236 17752 3292
rect 17752 3236 17756 3292
rect 17692 3232 17756 3236
rect 17772 3292 17836 3296
rect 17772 3236 17776 3292
rect 17776 3236 17832 3292
rect 17832 3236 17836 3292
rect 17772 3232 17836 3236
rect 17852 3292 17916 3296
rect 17852 3236 17856 3292
rect 17856 3236 17912 3292
rect 17912 3236 17916 3292
rect 17852 3232 17916 3236
rect 22612 3292 22676 3296
rect 22612 3236 22616 3292
rect 22616 3236 22672 3292
rect 22672 3236 22676 3292
rect 22612 3232 22676 3236
rect 22692 3292 22756 3296
rect 22692 3236 22696 3292
rect 22696 3236 22752 3292
rect 22752 3236 22756 3292
rect 22692 3232 22756 3236
rect 22772 3292 22836 3296
rect 22772 3236 22776 3292
rect 22776 3236 22832 3292
rect 22832 3236 22836 3292
rect 22772 3232 22836 3236
rect 22852 3292 22916 3296
rect 22852 3236 22856 3292
rect 22856 3236 22912 3292
rect 22912 3236 22916 3292
rect 22852 3232 22916 3236
rect 27612 3292 27676 3296
rect 27612 3236 27616 3292
rect 27616 3236 27672 3292
rect 27672 3236 27676 3292
rect 27612 3232 27676 3236
rect 27692 3292 27756 3296
rect 27692 3236 27696 3292
rect 27696 3236 27752 3292
rect 27752 3236 27756 3292
rect 27692 3232 27756 3236
rect 27772 3292 27836 3296
rect 27772 3236 27776 3292
rect 27776 3236 27832 3292
rect 27832 3236 27836 3292
rect 27772 3232 27836 3236
rect 27852 3292 27916 3296
rect 27852 3236 27856 3292
rect 27856 3236 27912 3292
rect 27912 3236 27916 3292
rect 27852 3232 27916 3236
rect 32612 3292 32676 3296
rect 32612 3236 32616 3292
rect 32616 3236 32672 3292
rect 32672 3236 32676 3292
rect 32612 3232 32676 3236
rect 32692 3292 32756 3296
rect 32692 3236 32696 3292
rect 32696 3236 32752 3292
rect 32752 3236 32756 3292
rect 32692 3232 32756 3236
rect 32772 3292 32836 3296
rect 32772 3236 32776 3292
rect 32776 3236 32832 3292
rect 32832 3236 32836 3292
rect 32772 3232 32836 3236
rect 32852 3292 32916 3296
rect 32852 3236 32856 3292
rect 32856 3236 32912 3292
rect 32912 3236 32916 3292
rect 32852 3232 32916 3236
rect 37612 3292 37676 3296
rect 37612 3236 37616 3292
rect 37616 3236 37672 3292
rect 37672 3236 37676 3292
rect 37612 3232 37676 3236
rect 37692 3292 37756 3296
rect 37692 3236 37696 3292
rect 37696 3236 37752 3292
rect 37752 3236 37756 3292
rect 37692 3232 37756 3236
rect 37772 3292 37836 3296
rect 37772 3236 37776 3292
rect 37776 3236 37832 3292
rect 37832 3236 37836 3292
rect 37772 3232 37836 3236
rect 37852 3292 37916 3296
rect 37852 3236 37856 3292
rect 37856 3236 37912 3292
rect 37912 3236 37916 3292
rect 37852 3232 37916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 6952 2748 7016 2752
rect 6952 2692 6956 2748
rect 6956 2692 7012 2748
rect 7012 2692 7016 2748
rect 6952 2688 7016 2692
rect 7032 2748 7096 2752
rect 7032 2692 7036 2748
rect 7036 2692 7092 2748
rect 7092 2692 7096 2748
rect 7032 2688 7096 2692
rect 7112 2748 7176 2752
rect 7112 2692 7116 2748
rect 7116 2692 7172 2748
rect 7172 2692 7176 2748
rect 7112 2688 7176 2692
rect 7192 2748 7256 2752
rect 7192 2692 7196 2748
rect 7196 2692 7252 2748
rect 7252 2692 7256 2748
rect 7192 2688 7256 2692
rect 11952 2748 12016 2752
rect 11952 2692 11956 2748
rect 11956 2692 12012 2748
rect 12012 2692 12016 2748
rect 11952 2688 12016 2692
rect 12032 2748 12096 2752
rect 12032 2692 12036 2748
rect 12036 2692 12092 2748
rect 12092 2692 12096 2748
rect 12032 2688 12096 2692
rect 12112 2748 12176 2752
rect 12112 2692 12116 2748
rect 12116 2692 12172 2748
rect 12172 2692 12176 2748
rect 12112 2688 12176 2692
rect 12192 2748 12256 2752
rect 12192 2692 12196 2748
rect 12196 2692 12252 2748
rect 12252 2692 12256 2748
rect 12192 2688 12256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 21952 2748 22016 2752
rect 21952 2692 21956 2748
rect 21956 2692 22012 2748
rect 22012 2692 22016 2748
rect 21952 2688 22016 2692
rect 22032 2748 22096 2752
rect 22032 2692 22036 2748
rect 22036 2692 22092 2748
rect 22092 2692 22096 2748
rect 22032 2688 22096 2692
rect 22112 2748 22176 2752
rect 22112 2692 22116 2748
rect 22116 2692 22172 2748
rect 22172 2692 22176 2748
rect 22112 2688 22176 2692
rect 22192 2748 22256 2752
rect 22192 2692 22196 2748
rect 22196 2692 22252 2748
rect 22252 2692 22256 2748
rect 22192 2688 22256 2692
rect 26952 2748 27016 2752
rect 26952 2692 26956 2748
rect 26956 2692 27012 2748
rect 27012 2692 27016 2748
rect 26952 2688 27016 2692
rect 27032 2748 27096 2752
rect 27032 2692 27036 2748
rect 27036 2692 27092 2748
rect 27092 2692 27096 2748
rect 27032 2688 27096 2692
rect 27112 2748 27176 2752
rect 27112 2692 27116 2748
rect 27116 2692 27172 2748
rect 27172 2692 27176 2748
rect 27112 2688 27176 2692
rect 27192 2748 27256 2752
rect 27192 2692 27196 2748
rect 27196 2692 27252 2748
rect 27252 2692 27256 2748
rect 27192 2688 27256 2692
rect 31952 2748 32016 2752
rect 31952 2692 31956 2748
rect 31956 2692 32012 2748
rect 32012 2692 32016 2748
rect 31952 2688 32016 2692
rect 32032 2748 32096 2752
rect 32032 2692 32036 2748
rect 32036 2692 32092 2748
rect 32092 2692 32096 2748
rect 32032 2688 32096 2692
rect 32112 2748 32176 2752
rect 32112 2692 32116 2748
rect 32116 2692 32172 2748
rect 32172 2692 32176 2748
rect 32112 2688 32176 2692
rect 32192 2748 32256 2752
rect 32192 2692 32196 2748
rect 32196 2692 32252 2748
rect 32252 2692 32256 2748
rect 32192 2688 32256 2692
rect 36952 2748 37016 2752
rect 36952 2692 36956 2748
rect 36956 2692 37012 2748
rect 37012 2692 37016 2748
rect 36952 2688 37016 2692
rect 37032 2748 37096 2752
rect 37032 2692 37036 2748
rect 37036 2692 37092 2748
rect 37092 2692 37096 2748
rect 37032 2688 37096 2692
rect 37112 2748 37176 2752
rect 37112 2692 37116 2748
rect 37116 2692 37172 2748
rect 37172 2692 37176 2748
rect 37112 2688 37176 2692
rect 37192 2748 37256 2752
rect 37192 2692 37196 2748
rect 37196 2692 37252 2748
rect 37252 2692 37256 2748
rect 37192 2688 37256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 7612 2204 7676 2208
rect 7612 2148 7616 2204
rect 7616 2148 7672 2204
rect 7672 2148 7676 2204
rect 7612 2144 7676 2148
rect 7692 2204 7756 2208
rect 7692 2148 7696 2204
rect 7696 2148 7752 2204
rect 7752 2148 7756 2204
rect 7692 2144 7756 2148
rect 7772 2204 7836 2208
rect 7772 2148 7776 2204
rect 7776 2148 7832 2204
rect 7832 2148 7836 2204
rect 7772 2144 7836 2148
rect 7852 2204 7916 2208
rect 7852 2148 7856 2204
rect 7856 2148 7912 2204
rect 7912 2148 7916 2204
rect 7852 2144 7916 2148
rect 12612 2204 12676 2208
rect 12612 2148 12616 2204
rect 12616 2148 12672 2204
rect 12672 2148 12676 2204
rect 12612 2144 12676 2148
rect 12692 2204 12756 2208
rect 12692 2148 12696 2204
rect 12696 2148 12752 2204
rect 12752 2148 12756 2204
rect 12692 2144 12756 2148
rect 12772 2204 12836 2208
rect 12772 2148 12776 2204
rect 12776 2148 12832 2204
rect 12832 2148 12836 2204
rect 12772 2144 12836 2148
rect 12852 2204 12916 2208
rect 12852 2148 12856 2204
rect 12856 2148 12912 2204
rect 12912 2148 12916 2204
rect 12852 2144 12916 2148
rect 17612 2204 17676 2208
rect 17612 2148 17616 2204
rect 17616 2148 17672 2204
rect 17672 2148 17676 2204
rect 17612 2144 17676 2148
rect 17692 2204 17756 2208
rect 17692 2148 17696 2204
rect 17696 2148 17752 2204
rect 17752 2148 17756 2204
rect 17692 2144 17756 2148
rect 17772 2204 17836 2208
rect 17772 2148 17776 2204
rect 17776 2148 17832 2204
rect 17832 2148 17836 2204
rect 17772 2144 17836 2148
rect 17852 2204 17916 2208
rect 17852 2148 17856 2204
rect 17856 2148 17912 2204
rect 17912 2148 17916 2204
rect 17852 2144 17916 2148
rect 22612 2204 22676 2208
rect 22612 2148 22616 2204
rect 22616 2148 22672 2204
rect 22672 2148 22676 2204
rect 22612 2144 22676 2148
rect 22692 2204 22756 2208
rect 22692 2148 22696 2204
rect 22696 2148 22752 2204
rect 22752 2148 22756 2204
rect 22692 2144 22756 2148
rect 22772 2204 22836 2208
rect 22772 2148 22776 2204
rect 22776 2148 22832 2204
rect 22832 2148 22836 2204
rect 22772 2144 22836 2148
rect 22852 2204 22916 2208
rect 22852 2148 22856 2204
rect 22856 2148 22912 2204
rect 22912 2148 22916 2204
rect 22852 2144 22916 2148
rect 27612 2204 27676 2208
rect 27612 2148 27616 2204
rect 27616 2148 27672 2204
rect 27672 2148 27676 2204
rect 27612 2144 27676 2148
rect 27692 2204 27756 2208
rect 27692 2148 27696 2204
rect 27696 2148 27752 2204
rect 27752 2148 27756 2204
rect 27692 2144 27756 2148
rect 27772 2204 27836 2208
rect 27772 2148 27776 2204
rect 27776 2148 27832 2204
rect 27832 2148 27836 2204
rect 27772 2144 27836 2148
rect 27852 2204 27916 2208
rect 27852 2148 27856 2204
rect 27856 2148 27912 2204
rect 27912 2148 27916 2204
rect 27852 2144 27916 2148
rect 32612 2204 32676 2208
rect 32612 2148 32616 2204
rect 32616 2148 32672 2204
rect 32672 2148 32676 2204
rect 32612 2144 32676 2148
rect 32692 2204 32756 2208
rect 32692 2148 32696 2204
rect 32696 2148 32752 2204
rect 32752 2148 32756 2204
rect 32692 2144 32756 2148
rect 32772 2204 32836 2208
rect 32772 2148 32776 2204
rect 32776 2148 32832 2204
rect 32832 2148 32836 2204
rect 32772 2144 32836 2148
rect 32852 2204 32916 2208
rect 32852 2148 32856 2204
rect 32856 2148 32912 2204
rect 32912 2148 32916 2204
rect 32852 2144 32916 2148
rect 37612 2204 37676 2208
rect 37612 2148 37616 2204
rect 37616 2148 37672 2204
rect 37672 2148 37676 2204
rect 37612 2144 37676 2148
rect 37692 2204 37756 2208
rect 37692 2148 37696 2204
rect 37696 2148 37752 2204
rect 37752 2148 37756 2204
rect 37692 2144 37756 2148
rect 37772 2204 37836 2208
rect 37772 2148 37776 2204
rect 37776 2148 37832 2204
rect 37832 2148 37836 2204
rect 37772 2144 37836 2148
rect 37852 2204 37916 2208
rect 37852 2148 37856 2204
rect 37856 2148 37912 2204
rect 37912 2148 37916 2204
rect 37852 2144 37916 2148
<< metal4 >>
rect 1944 37568 2264 37584
rect 1944 37504 1952 37568
rect 2016 37504 2032 37568
rect 2096 37504 2112 37568
rect 2176 37504 2192 37568
rect 2256 37504 2264 37568
rect 1944 36480 2264 37504
rect 1944 36416 1952 36480
rect 2016 36416 2032 36480
rect 2096 36416 2112 36480
rect 2176 36416 2192 36480
rect 2256 36416 2264 36480
rect 1944 35392 2264 36416
rect 1944 35328 1952 35392
rect 2016 35328 2032 35392
rect 2096 35328 2112 35392
rect 2176 35328 2192 35392
rect 2256 35328 2264 35392
rect 1944 34304 2264 35328
rect 1944 34240 1952 34304
rect 2016 34240 2032 34304
rect 2096 34240 2112 34304
rect 2176 34240 2192 34304
rect 2256 34240 2264 34304
rect 1944 33294 2264 34240
rect 1944 33216 1986 33294
rect 2222 33216 2264 33294
rect 1944 33152 1952 33216
rect 2256 33152 2264 33216
rect 1944 33058 1986 33152
rect 2222 33058 2264 33152
rect 1944 32128 2264 33058
rect 1944 32064 1952 32128
rect 2016 32064 2032 32128
rect 2096 32064 2112 32128
rect 2176 32064 2192 32128
rect 2256 32064 2264 32128
rect 1944 31040 2264 32064
rect 1944 30976 1952 31040
rect 2016 30976 2032 31040
rect 2096 30976 2112 31040
rect 2176 30976 2192 31040
rect 2256 30976 2264 31040
rect 1944 29952 2264 30976
rect 1944 29888 1952 29952
rect 2016 29888 2032 29952
rect 2096 29888 2112 29952
rect 2176 29888 2192 29952
rect 2256 29888 2264 29952
rect 1944 28864 2264 29888
rect 1944 28800 1952 28864
rect 2016 28800 2032 28864
rect 2096 28800 2112 28864
rect 2176 28800 2192 28864
rect 2256 28800 2264 28864
rect 1944 28294 2264 28800
rect 1944 28058 1986 28294
rect 2222 28058 2264 28294
rect 1944 27776 2264 28058
rect 1944 27712 1952 27776
rect 2016 27712 2032 27776
rect 2096 27712 2112 27776
rect 2176 27712 2192 27776
rect 2256 27712 2264 27776
rect 1944 26688 2264 27712
rect 1944 26624 1952 26688
rect 2016 26624 2032 26688
rect 2096 26624 2112 26688
rect 2176 26624 2192 26688
rect 2256 26624 2264 26688
rect 1944 25600 2264 26624
rect 1944 25536 1952 25600
rect 2016 25536 2032 25600
rect 2096 25536 2112 25600
rect 2176 25536 2192 25600
rect 2256 25536 2264 25600
rect 1944 24512 2264 25536
rect 1944 24448 1952 24512
rect 2016 24448 2032 24512
rect 2096 24448 2112 24512
rect 2176 24448 2192 24512
rect 2256 24448 2264 24512
rect 1944 23424 2264 24448
rect 1944 23360 1952 23424
rect 2016 23360 2032 23424
rect 2096 23360 2112 23424
rect 2176 23360 2192 23424
rect 2256 23360 2264 23424
rect 1944 23294 2264 23360
rect 1944 23058 1986 23294
rect 2222 23058 2264 23294
rect 1944 22336 2264 23058
rect 1944 22272 1952 22336
rect 2016 22272 2032 22336
rect 2096 22272 2112 22336
rect 2176 22272 2192 22336
rect 2256 22272 2264 22336
rect 1944 21248 2264 22272
rect 1944 21184 1952 21248
rect 2016 21184 2032 21248
rect 2096 21184 2112 21248
rect 2176 21184 2192 21248
rect 2256 21184 2264 21248
rect 1944 20160 2264 21184
rect 1944 20096 1952 20160
rect 2016 20096 2032 20160
rect 2096 20096 2112 20160
rect 2176 20096 2192 20160
rect 2256 20096 2264 20160
rect 1944 19072 2264 20096
rect 1944 19008 1952 19072
rect 2016 19008 2032 19072
rect 2096 19008 2112 19072
rect 2176 19008 2192 19072
rect 2256 19008 2264 19072
rect 1944 18294 2264 19008
rect 1944 18058 1986 18294
rect 2222 18058 2264 18294
rect 1944 17984 2264 18058
rect 1944 17920 1952 17984
rect 2016 17920 2032 17984
rect 2096 17920 2112 17984
rect 2176 17920 2192 17984
rect 2256 17920 2264 17984
rect 1944 16896 2264 17920
rect 1944 16832 1952 16896
rect 2016 16832 2032 16896
rect 2096 16832 2112 16896
rect 2176 16832 2192 16896
rect 2256 16832 2264 16896
rect 1944 15808 2264 16832
rect 1944 15744 1952 15808
rect 2016 15744 2032 15808
rect 2096 15744 2112 15808
rect 2176 15744 2192 15808
rect 2256 15744 2264 15808
rect 1944 14720 2264 15744
rect 1944 14656 1952 14720
rect 2016 14656 2032 14720
rect 2096 14656 2112 14720
rect 2176 14656 2192 14720
rect 2256 14656 2264 14720
rect 1944 13632 2264 14656
rect 1944 13568 1952 13632
rect 2016 13568 2032 13632
rect 2096 13568 2112 13632
rect 2176 13568 2192 13632
rect 2256 13568 2264 13632
rect 1944 13294 2264 13568
rect 1944 13058 1986 13294
rect 2222 13058 2264 13294
rect 1944 12544 2264 13058
rect 1944 12480 1952 12544
rect 2016 12480 2032 12544
rect 2096 12480 2112 12544
rect 2176 12480 2192 12544
rect 2256 12480 2264 12544
rect 1944 11456 2264 12480
rect 1944 11392 1952 11456
rect 2016 11392 2032 11456
rect 2096 11392 2112 11456
rect 2176 11392 2192 11456
rect 2256 11392 2264 11456
rect 1944 10368 2264 11392
rect 1944 10304 1952 10368
rect 2016 10304 2032 10368
rect 2096 10304 2112 10368
rect 2176 10304 2192 10368
rect 2256 10304 2264 10368
rect 1944 9280 2264 10304
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8294 2264 9216
rect 1944 8192 1986 8294
rect 2222 8192 2264 8294
rect 1944 8128 1952 8192
rect 2256 8128 2264 8192
rect 1944 8058 1986 8128
rect 2222 8058 2264 8128
rect 1944 7104 2264 8058
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3294 2264 3776
rect 1944 3058 1986 3294
rect 2222 3058 2264 3294
rect 1944 2752 2264 3058
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 37024 2924 37584
rect 2604 36960 2612 37024
rect 2676 36960 2692 37024
rect 2756 36960 2772 37024
rect 2836 36960 2852 37024
rect 2916 36960 2924 37024
rect 2604 35936 2924 36960
rect 2604 35872 2612 35936
rect 2676 35872 2692 35936
rect 2756 35872 2772 35936
rect 2836 35872 2852 35936
rect 2916 35872 2924 35936
rect 2604 34848 2924 35872
rect 2604 34784 2612 34848
rect 2676 34784 2692 34848
rect 2756 34784 2772 34848
rect 2836 34784 2852 34848
rect 2916 34784 2924 34848
rect 2604 33954 2924 34784
rect 2604 33760 2646 33954
rect 2882 33760 2924 33954
rect 2604 33696 2612 33760
rect 2676 33696 2692 33718
rect 2756 33696 2772 33718
rect 2836 33696 2852 33718
rect 2916 33696 2924 33760
rect 2604 32672 2924 33696
rect 2604 32608 2612 32672
rect 2676 32608 2692 32672
rect 2756 32608 2772 32672
rect 2836 32608 2852 32672
rect 2916 32608 2924 32672
rect 2604 31584 2924 32608
rect 2604 31520 2612 31584
rect 2676 31520 2692 31584
rect 2756 31520 2772 31584
rect 2836 31520 2852 31584
rect 2916 31520 2924 31584
rect 2604 30496 2924 31520
rect 2604 30432 2612 30496
rect 2676 30432 2692 30496
rect 2756 30432 2772 30496
rect 2836 30432 2852 30496
rect 2916 30432 2924 30496
rect 2604 29408 2924 30432
rect 2604 29344 2612 29408
rect 2676 29344 2692 29408
rect 2756 29344 2772 29408
rect 2836 29344 2852 29408
rect 2916 29344 2924 29408
rect 2604 28954 2924 29344
rect 2604 28718 2646 28954
rect 2882 28718 2924 28954
rect 2604 28320 2924 28718
rect 2604 28256 2612 28320
rect 2676 28256 2692 28320
rect 2756 28256 2772 28320
rect 2836 28256 2852 28320
rect 2916 28256 2924 28320
rect 2604 27232 2924 28256
rect 2604 27168 2612 27232
rect 2676 27168 2692 27232
rect 2756 27168 2772 27232
rect 2836 27168 2852 27232
rect 2916 27168 2924 27232
rect 2604 26144 2924 27168
rect 2604 26080 2612 26144
rect 2676 26080 2692 26144
rect 2756 26080 2772 26144
rect 2836 26080 2852 26144
rect 2916 26080 2924 26144
rect 2604 25056 2924 26080
rect 2604 24992 2612 25056
rect 2676 24992 2692 25056
rect 2756 24992 2772 25056
rect 2836 24992 2852 25056
rect 2916 24992 2924 25056
rect 2604 23968 2924 24992
rect 2604 23904 2612 23968
rect 2676 23954 2692 23968
rect 2756 23954 2772 23968
rect 2836 23954 2852 23968
rect 2916 23904 2924 23968
rect 2604 23718 2646 23904
rect 2882 23718 2924 23904
rect 2604 22880 2924 23718
rect 2604 22816 2612 22880
rect 2676 22816 2692 22880
rect 2756 22816 2772 22880
rect 2836 22816 2852 22880
rect 2916 22816 2924 22880
rect 2604 21792 2924 22816
rect 2604 21728 2612 21792
rect 2676 21728 2692 21792
rect 2756 21728 2772 21792
rect 2836 21728 2852 21792
rect 2916 21728 2924 21792
rect 2604 20704 2924 21728
rect 2604 20640 2612 20704
rect 2676 20640 2692 20704
rect 2756 20640 2772 20704
rect 2836 20640 2852 20704
rect 2916 20640 2924 20704
rect 2604 19616 2924 20640
rect 2604 19552 2612 19616
rect 2676 19552 2692 19616
rect 2756 19552 2772 19616
rect 2836 19552 2852 19616
rect 2916 19552 2924 19616
rect 2604 18954 2924 19552
rect 2604 18718 2646 18954
rect 2882 18718 2924 18954
rect 2604 18528 2924 18718
rect 2604 18464 2612 18528
rect 2676 18464 2692 18528
rect 2756 18464 2772 18528
rect 2836 18464 2852 18528
rect 2916 18464 2924 18528
rect 2604 17440 2924 18464
rect 2604 17376 2612 17440
rect 2676 17376 2692 17440
rect 2756 17376 2772 17440
rect 2836 17376 2852 17440
rect 2916 17376 2924 17440
rect 2604 16352 2924 17376
rect 2604 16288 2612 16352
rect 2676 16288 2692 16352
rect 2756 16288 2772 16352
rect 2836 16288 2852 16352
rect 2916 16288 2924 16352
rect 2604 15264 2924 16288
rect 2604 15200 2612 15264
rect 2676 15200 2692 15264
rect 2756 15200 2772 15264
rect 2836 15200 2852 15264
rect 2916 15200 2924 15264
rect 2604 14176 2924 15200
rect 2604 14112 2612 14176
rect 2676 14112 2692 14176
rect 2756 14112 2772 14176
rect 2836 14112 2852 14176
rect 2916 14112 2924 14176
rect 2604 13954 2924 14112
rect 2604 13718 2646 13954
rect 2882 13718 2924 13954
rect 2604 13088 2924 13718
rect 2604 13024 2612 13088
rect 2676 13024 2692 13088
rect 2756 13024 2772 13088
rect 2836 13024 2852 13088
rect 2916 13024 2924 13088
rect 2604 12000 2924 13024
rect 2604 11936 2612 12000
rect 2676 11936 2692 12000
rect 2756 11936 2772 12000
rect 2836 11936 2852 12000
rect 2916 11936 2924 12000
rect 2604 10912 2924 11936
rect 2604 10848 2612 10912
rect 2676 10848 2692 10912
rect 2756 10848 2772 10912
rect 2836 10848 2852 10912
rect 2916 10848 2924 10912
rect 2604 9824 2924 10848
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 8954 2924 9760
rect 2604 8736 2646 8954
rect 2882 8736 2924 8954
rect 2604 8672 2612 8736
rect 2676 8672 2692 8718
rect 2756 8672 2772 8718
rect 2836 8672 2852 8718
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3954 2924 4320
rect 2604 3718 2646 3954
rect 2882 3718 2924 3954
rect 2604 3296 2924 3718
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 6944 37568 7264 37584
rect 6944 37504 6952 37568
rect 7016 37504 7032 37568
rect 7096 37504 7112 37568
rect 7176 37504 7192 37568
rect 7256 37504 7264 37568
rect 6944 36480 7264 37504
rect 6944 36416 6952 36480
rect 7016 36416 7032 36480
rect 7096 36416 7112 36480
rect 7176 36416 7192 36480
rect 7256 36416 7264 36480
rect 6944 35392 7264 36416
rect 6944 35328 6952 35392
rect 7016 35328 7032 35392
rect 7096 35328 7112 35392
rect 7176 35328 7192 35392
rect 7256 35328 7264 35392
rect 6944 34304 7264 35328
rect 6944 34240 6952 34304
rect 7016 34240 7032 34304
rect 7096 34240 7112 34304
rect 7176 34240 7192 34304
rect 7256 34240 7264 34304
rect 6944 33294 7264 34240
rect 6944 33216 6986 33294
rect 7222 33216 7264 33294
rect 6944 33152 6952 33216
rect 7256 33152 7264 33216
rect 6944 33058 6986 33152
rect 7222 33058 7264 33152
rect 6944 32128 7264 33058
rect 6944 32064 6952 32128
rect 7016 32064 7032 32128
rect 7096 32064 7112 32128
rect 7176 32064 7192 32128
rect 7256 32064 7264 32128
rect 6944 31040 7264 32064
rect 6944 30976 6952 31040
rect 7016 30976 7032 31040
rect 7096 30976 7112 31040
rect 7176 30976 7192 31040
rect 7256 30976 7264 31040
rect 6944 29952 7264 30976
rect 6944 29888 6952 29952
rect 7016 29888 7032 29952
rect 7096 29888 7112 29952
rect 7176 29888 7192 29952
rect 7256 29888 7264 29952
rect 6944 28864 7264 29888
rect 6944 28800 6952 28864
rect 7016 28800 7032 28864
rect 7096 28800 7112 28864
rect 7176 28800 7192 28864
rect 7256 28800 7264 28864
rect 6944 28294 7264 28800
rect 6944 28058 6986 28294
rect 7222 28058 7264 28294
rect 6944 27776 7264 28058
rect 6944 27712 6952 27776
rect 7016 27712 7032 27776
rect 7096 27712 7112 27776
rect 7176 27712 7192 27776
rect 7256 27712 7264 27776
rect 6944 26688 7264 27712
rect 6944 26624 6952 26688
rect 7016 26624 7032 26688
rect 7096 26624 7112 26688
rect 7176 26624 7192 26688
rect 7256 26624 7264 26688
rect 6944 25600 7264 26624
rect 6944 25536 6952 25600
rect 7016 25536 7032 25600
rect 7096 25536 7112 25600
rect 7176 25536 7192 25600
rect 7256 25536 7264 25600
rect 6944 24512 7264 25536
rect 6944 24448 6952 24512
rect 7016 24448 7032 24512
rect 7096 24448 7112 24512
rect 7176 24448 7192 24512
rect 7256 24448 7264 24512
rect 6944 23424 7264 24448
rect 6944 23360 6952 23424
rect 7016 23360 7032 23424
rect 7096 23360 7112 23424
rect 7176 23360 7192 23424
rect 7256 23360 7264 23424
rect 6944 23294 7264 23360
rect 6944 23058 6986 23294
rect 7222 23058 7264 23294
rect 6944 22336 7264 23058
rect 6944 22272 6952 22336
rect 7016 22272 7032 22336
rect 7096 22272 7112 22336
rect 7176 22272 7192 22336
rect 7256 22272 7264 22336
rect 6944 21248 7264 22272
rect 6944 21184 6952 21248
rect 7016 21184 7032 21248
rect 7096 21184 7112 21248
rect 7176 21184 7192 21248
rect 7256 21184 7264 21248
rect 6944 20160 7264 21184
rect 6944 20096 6952 20160
rect 7016 20096 7032 20160
rect 7096 20096 7112 20160
rect 7176 20096 7192 20160
rect 7256 20096 7264 20160
rect 6944 19072 7264 20096
rect 6944 19008 6952 19072
rect 7016 19008 7032 19072
rect 7096 19008 7112 19072
rect 7176 19008 7192 19072
rect 7256 19008 7264 19072
rect 6944 18294 7264 19008
rect 6944 18058 6986 18294
rect 7222 18058 7264 18294
rect 6944 17984 7264 18058
rect 6944 17920 6952 17984
rect 7016 17920 7032 17984
rect 7096 17920 7112 17984
rect 7176 17920 7192 17984
rect 7256 17920 7264 17984
rect 6944 16896 7264 17920
rect 6944 16832 6952 16896
rect 7016 16832 7032 16896
rect 7096 16832 7112 16896
rect 7176 16832 7192 16896
rect 7256 16832 7264 16896
rect 6944 15808 7264 16832
rect 6944 15744 6952 15808
rect 7016 15744 7032 15808
rect 7096 15744 7112 15808
rect 7176 15744 7192 15808
rect 7256 15744 7264 15808
rect 6944 14720 7264 15744
rect 6944 14656 6952 14720
rect 7016 14656 7032 14720
rect 7096 14656 7112 14720
rect 7176 14656 7192 14720
rect 7256 14656 7264 14720
rect 6944 13632 7264 14656
rect 6944 13568 6952 13632
rect 7016 13568 7032 13632
rect 7096 13568 7112 13632
rect 7176 13568 7192 13632
rect 7256 13568 7264 13632
rect 6944 13294 7264 13568
rect 6944 13058 6986 13294
rect 7222 13058 7264 13294
rect 6944 12544 7264 13058
rect 6944 12480 6952 12544
rect 7016 12480 7032 12544
rect 7096 12480 7112 12544
rect 7176 12480 7192 12544
rect 7256 12480 7264 12544
rect 6944 11456 7264 12480
rect 6944 11392 6952 11456
rect 7016 11392 7032 11456
rect 7096 11392 7112 11456
rect 7176 11392 7192 11456
rect 7256 11392 7264 11456
rect 6944 10368 7264 11392
rect 6944 10304 6952 10368
rect 7016 10304 7032 10368
rect 7096 10304 7112 10368
rect 7176 10304 7192 10368
rect 7256 10304 7264 10368
rect 6944 9280 7264 10304
rect 6944 9216 6952 9280
rect 7016 9216 7032 9280
rect 7096 9216 7112 9280
rect 7176 9216 7192 9280
rect 7256 9216 7264 9280
rect 6944 8294 7264 9216
rect 6944 8192 6986 8294
rect 7222 8192 7264 8294
rect 6944 8128 6952 8192
rect 7256 8128 7264 8192
rect 6944 8058 6986 8128
rect 7222 8058 7264 8128
rect 6944 7104 7264 8058
rect 6944 7040 6952 7104
rect 7016 7040 7032 7104
rect 7096 7040 7112 7104
rect 7176 7040 7192 7104
rect 7256 7040 7264 7104
rect 6944 6016 7264 7040
rect 6944 5952 6952 6016
rect 7016 5952 7032 6016
rect 7096 5952 7112 6016
rect 7176 5952 7192 6016
rect 7256 5952 7264 6016
rect 6944 4928 7264 5952
rect 6944 4864 6952 4928
rect 7016 4864 7032 4928
rect 7096 4864 7112 4928
rect 7176 4864 7192 4928
rect 7256 4864 7264 4928
rect 6944 3840 7264 4864
rect 6944 3776 6952 3840
rect 7016 3776 7032 3840
rect 7096 3776 7112 3840
rect 7176 3776 7192 3840
rect 7256 3776 7264 3840
rect 6944 3294 7264 3776
rect 6944 3058 6986 3294
rect 7222 3058 7264 3294
rect 6944 2752 7264 3058
rect 6944 2688 6952 2752
rect 7016 2688 7032 2752
rect 7096 2688 7112 2752
rect 7176 2688 7192 2752
rect 7256 2688 7264 2752
rect 6944 2128 7264 2688
rect 7604 37024 7924 37584
rect 7604 36960 7612 37024
rect 7676 36960 7692 37024
rect 7756 36960 7772 37024
rect 7836 36960 7852 37024
rect 7916 36960 7924 37024
rect 7604 35936 7924 36960
rect 7604 35872 7612 35936
rect 7676 35872 7692 35936
rect 7756 35872 7772 35936
rect 7836 35872 7852 35936
rect 7916 35872 7924 35936
rect 7604 34848 7924 35872
rect 7604 34784 7612 34848
rect 7676 34784 7692 34848
rect 7756 34784 7772 34848
rect 7836 34784 7852 34848
rect 7916 34784 7924 34848
rect 7604 33954 7924 34784
rect 7604 33760 7646 33954
rect 7882 33760 7924 33954
rect 7604 33696 7612 33760
rect 7676 33696 7692 33718
rect 7756 33696 7772 33718
rect 7836 33696 7852 33718
rect 7916 33696 7924 33760
rect 7604 32672 7924 33696
rect 7604 32608 7612 32672
rect 7676 32608 7692 32672
rect 7756 32608 7772 32672
rect 7836 32608 7852 32672
rect 7916 32608 7924 32672
rect 7604 31584 7924 32608
rect 7604 31520 7612 31584
rect 7676 31520 7692 31584
rect 7756 31520 7772 31584
rect 7836 31520 7852 31584
rect 7916 31520 7924 31584
rect 7604 30496 7924 31520
rect 7604 30432 7612 30496
rect 7676 30432 7692 30496
rect 7756 30432 7772 30496
rect 7836 30432 7852 30496
rect 7916 30432 7924 30496
rect 7604 29408 7924 30432
rect 7604 29344 7612 29408
rect 7676 29344 7692 29408
rect 7756 29344 7772 29408
rect 7836 29344 7852 29408
rect 7916 29344 7924 29408
rect 7604 28954 7924 29344
rect 7604 28718 7646 28954
rect 7882 28718 7924 28954
rect 7604 28320 7924 28718
rect 7604 28256 7612 28320
rect 7676 28256 7692 28320
rect 7756 28256 7772 28320
rect 7836 28256 7852 28320
rect 7916 28256 7924 28320
rect 7604 27232 7924 28256
rect 7604 27168 7612 27232
rect 7676 27168 7692 27232
rect 7756 27168 7772 27232
rect 7836 27168 7852 27232
rect 7916 27168 7924 27232
rect 7604 26144 7924 27168
rect 7604 26080 7612 26144
rect 7676 26080 7692 26144
rect 7756 26080 7772 26144
rect 7836 26080 7852 26144
rect 7916 26080 7924 26144
rect 7604 25056 7924 26080
rect 7604 24992 7612 25056
rect 7676 24992 7692 25056
rect 7756 24992 7772 25056
rect 7836 24992 7852 25056
rect 7916 24992 7924 25056
rect 7604 23968 7924 24992
rect 7604 23904 7612 23968
rect 7676 23954 7692 23968
rect 7756 23954 7772 23968
rect 7836 23954 7852 23968
rect 7916 23904 7924 23968
rect 7604 23718 7646 23904
rect 7882 23718 7924 23904
rect 7604 22880 7924 23718
rect 7604 22816 7612 22880
rect 7676 22816 7692 22880
rect 7756 22816 7772 22880
rect 7836 22816 7852 22880
rect 7916 22816 7924 22880
rect 7604 21792 7924 22816
rect 7604 21728 7612 21792
rect 7676 21728 7692 21792
rect 7756 21728 7772 21792
rect 7836 21728 7852 21792
rect 7916 21728 7924 21792
rect 7604 20704 7924 21728
rect 7604 20640 7612 20704
rect 7676 20640 7692 20704
rect 7756 20640 7772 20704
rect 7836 20640 7852 20704
rect 7916 20640 7924 20704
rect 7604 19616 7924 20640
rect 7604 19552 7612 19616
rect 7676 19552 7692 19616
rect 7756 19552 7772 19616
rect 7836 19552 7852 19616
rect 7916 19552 7924 19616
rect 7604 18954 7924 19552
rect 7604 18718 7646 18954
rect 7882 18718 7924 18954
rect 7604 18528 7924 18718
rect 7604 18464 7612 18528
rect 7676 18464 7692 18528
rect 7756 18464 7772 18528
rect 7836 18464 7852 18528
rect 7916 18464 7924 18528
rect 7604 17440 7924 18464
rect 7604 17376 7612 17440
rect 7676 17376 7692 17440
rect 7756 17376 7772 17440
rect 7836 17376 7852 17440
rect 7916 17376 7924 17440
rect 7604 16352 7924 17376
rect 7604 16288 7612 16352
rect 7676 16288 7692 16352
rect 7756 16288 7772 16352
rect 7836 16288 7852 16352
rect 7916 16288 7924 16352
rect 7604 15264 7924 16288
rect 7604 15200 7612 15264
rect 7676 15200 7692 15264
rect 7756 15200 7772 15264
rect 7836 15200 7852 15264
rect 7916 15200 7924 15264
rect 7604 14176 7924 15200
rect 7604 14112 7612 14176
rect 7676 14112 7692 14176
rect 7756 14112 7772 14176
rect 7836 14112 7852 14176
rect 7916 14112 7924 14176
rect 7604 13954 7924 14112
rect 7604 13718 7646 13954
rect 7882 13718 7924 13954
rect 7604 13088 7924 13718
rect 7604 13024 7612 13088
rect 7676 13024 7692 13088
rect 7756 13024 7772 13088
rect 7836 13024 7852 13088
rect 7916 13024 7924 13088
rect 7604 12000 7924 13024
rect 7604 11936 7612 12000
rect 7676 11936 7692 12000
rect 7756 11936 7772 12000
rect 7836 11936 7852 12000
rect 7916 11936 7924 12000
rect 7604 10912 7924 11936
rect 7604 10848 7612 10912
rect 7676 10848 7692 10912
rect 7756 10848 7772 10912
rect 7836 10848 7852 10912
rect 7916 10848 7924 10912
rect 7604 9824 7924 10848
rect 7604 9760 7612 9824
rect 7676 9760 7692 9824
rect 7756 9760 7772 9824
rect 7836 9760 7852 9824
rect 7916 9760 7924 9824
rect 7604 8954 7924 9760
rect 7604 8736 7646 8954
rect 7882 8736 7924 8954
rect 7604 8672 7612 8736
rect 7676 8672 7692 8718
rect 7756 8672 7772 8718
rect 7836 8672 7852 8718
rect 7916 8672 7924 8736
rect 7604 7648 7924 8672
rect 7604 7584 7612 7648
rect 7676 7584 7692 7648
rect 7756 7584 7772 7648
rect 7836 7584 7852 7648
rect 7916 7584 7924 7648
rect 7604 6560 7924 7584
rect 7604 6496 7612 6560
rect 7676 6496 7692 6560
rect 7756 6496 7772 6560
rect 7836 6496 7852 6560
rect 7916 6496 7924 6560
rect 7604 5472 7924 6496
rect 7604 5408 7612 5472
rect 7676 5408 7692 5472
rect 7756 5408 7772 5472
rect 7836 5408 7852 5472
rect 7916 5408 7924 5472
rect 7604 4384 7924 5408
rect 7604 4320 7612 4384
rect 7676 4320 7692 4384
rect 7756 4320 7772 4384
rect 7836 4320 7852 4384
rect 7916 4320 7924 4384
rect 7604 3954 7924 4320
rect 7604 3718 7646 3954
rect 7882 3718 7924 3954
rect 7604 3296 7924 3718
rect 7604 3232 7612 3296
rect 7676 3232 7692 3296
rect 7756 3232 7772 3296
rect 7836 3232 7852 3296
rect 7916 3232 7924 3296
rect 7604 2208 7924 3232
rect 7604 2144 7612 2208
rect 7676 2144 7692 2208
rect 7756 2144 7772 2208
rect 7836 2144 7852 2208
rect 7916 2144 7924 2208
rect 7604 2128 7924 2144
rect 11944 37568 12264 37584
rect 11944 37504 11952 37568
rect 12016 37504 12032 37568
rect 12096 37504 12112 37568
rect 12176 37504 12192 37568
rect 12256 37504 12264 37568
rect 11944 36480 12264 37504
rect 11944 36416 11952 36480
rect 12016 36416 12032 36480
rect 12096 36416 12112 36480
rect 12176 36416 12192 36480
rect 12256 36416 12264 36480
rect 11944 35392 12264 36416
rect 11944 35328 11952 35392
rect 12016 35328 12032 35392
rect 12096 35328 12112 35392
rect 12176 35328 12192 35392
rect 12256 35328 12264 35392
rect 11944 34304 12264 35328
rect 11944 34240 11952 34304
rect 12016 34240 12032 34304
rect 12096 34240 12112 34304
rect 12176 34240 12192 34304
rect 12256 34240 12264 34304
rect 11944 33294 12264 34240
rect 11944 33216 11986 33294
rect 12222 33216 12264 33294
rect 11944 33152 11952 33216
rect 12256 33152 12264 33216
rect 11944 33058 11986 33152
rect 12222 33058 12264 33152
rect 11944 32128 12264 33058
rect 11944 32064 11952 32128
rect 12016 32064 12032 32128
rect 12096 32064 12112 32128
rect 12176 32064 12192 32128
rect 12256 32064 12264 32128
rect 11944 31040 12264 32064
rect 11944 30976 11952 31040
rect 12016 30976 12032 31040
rect 12096 30976 12112 31040
rect 12176 30976 12192 31040
rect 12256 30976 12264 31040
rect 11944 29952 12264 30976
rect 11944 29888 11952 29952
rect 12016 29888 12032 29952
rect 12096 29888 12112 29952
rect 12176 29888 12192 29952
rect 12256 29888 12264 29952
rect 11944 28864 12264 29888
rect 11944 28800 11952 28864
rect 12016 28800 12032 28864
rect 12096 28800 12112 28864
rect 12176 28800 12192 28864
rect 12256 28800 12264 28864
rect 11944 28294 12264 28800
rect 11944 28058 11986 28294
rect 12222 28058 12264 28294
rect 11944 27776 12264 28058
rect 11944 27712 11952 27776
rect 12016 27712 12032 27776
rect 12096 27712 12112 27776
rect 12176 27712 12192 27776
rect 12256 27712 12264 27776
rect 11944 26688 12264 27712
rect 11944 26624 11952 26688
rect 12016 26624 12032 26688
rect 12096 26624 12112 26688
rect 12176 26624 12192 26688
rect 12256 26624 12264 26688
rect 11944 25600 12264 26624
rect 11944 25536 11952 25600
rect 12016 25536 12032 25600
rect 12096 25536 12112 25600
rect 12176 25536 12192 25600
rect 12256 25536 12264 25600
rect 11944 24512 12264 25536
rect 11944 24448 11952 24512
rect 12016 24448 12032 24512
rect 12096 24448 12112 24512
rect 12176 24448 12192 24512
rect 12256 24448 12264 24512
rect 11944 23424 12264 24448
rect 11944 23360 11952 23424
rect 12016 23360 12032 23424
rect 12096 23360 12112 23424
rect 12176 23360 12192 23424
rect 12256 23360 12264 23424
rect 11944 23294 12264 23360
rect 11944 23058 11986 23294
rect 12222 23058 12264 23294
rect 11944 22336 12264 23058
rect 11944 22272 11952 22336
rect 12016 22272 12032 22336
rect 12096 22272 12112 22336
rect 12176 22272 12192 22336
rect 12256 22272 12264 22336
rect 11944 21248 12264 22272
rect 11944 21184 11952 21248
rect 12016 21184 12032 21248
rect 12096 21184 12112 21248
rect 12176 21184 12192 21248
rect 12256 21184 12264 21248
rect 11944 20160 12264 21184
rect 11944 20096 11952 20160
rect 12016 20096 12032 20160
rect 12096 20096 12112 20160
rect 12176 20096 12192 20160
rect 12256 20096 12264 20160
rect 11944 19072 12264 20096
rect 11944 19008 11952 19072
rect 12016 19008 12032 19072
rect 12096 19008 12112 19072
rect 12176 19008 12192 19072
rect 12256 19008 12264 19072
rect 11944 18294 12264 19008
rect 11944 18058 11986 18294
rect 12222 18058 12264 18294
rect 11944 17984 12264 18058
rect 11944 17920 11952 17984
rect 12016 17920 12032 17984
rect 12096 17920 12112 17984
rect 12176 17920 12192 17984
rect 12256 17920 12264 17984
rect 11944 16896 12264 17920
rect 11944 16832 11952 16896
rect 12016 16832 12032 16896
rect 12096 16832 12112 16896
rect 12176 16832 12192 16896
rect 12256 16832 12264 16896
rect 11944 15808 12264 16832
rect 11944 15744 11952 15808
rect 12016 15744 12032 15808
rect 12096 15744 12112 15808
rect 12176 15744 12192 15808
rect 12256 15744 12264 15808
rect 11944 14720 12264 15744
rect 11944 14656 11952 14720
rect 12016 14656 12032 14720
rect 12096 14656 12112 14720
rect 12176 14656 12192 14720
rect 12256 14656 12264 14720
rect 11944 13632 12264 14656
rect 11944 13568 11952 13632
rect 12016 13568 12032 13632
rect 12096 13568 12112 13632
rect 12176 13568 12192 13632
rect 12256 13568 12264 13632
rect 11944 13294 12264 13568
rect 11944 13058 11986 13294
rect 12222 13058 12264 13294
rect 11944 12544 12264 13058
rect 11944 12480 11952 12544
rect 12016 12480 12032 12544
rect 12096 12480 12112 12544
rect 12176 12480 12192 12544
rect 12256 12480 12264 12544
rect 11944 11456 12264 12480
rect 11944 11392 11952 11456
rect 12016 11392 12032 11456
rect 12096 11392 12112 11456
rect 12176 11392 12192 11456
rect 12256 11392 12264 11456
rect 11944 10368 12264 11392
rect 11944 10304 11952 10368
rect 12016 10304 12032 10368
rect 12096 10304 12112 10368
rect 12176 10304 12192 10368
rect 12256 10304 12264 10368
rect 11944 9280 12264 10304
rect 11944 9216 11952 9280
rect 12016 9216 12032 9280
rect 12096 9216 12112 9280
rect 12176 9216 12192 9280
rect 12256 9216 12264 9280
rect 11944 8294 12264 9216
rect 11944 8192 11986 8294
rect 12222 8192 12264 8294
rect 11944 8128 11952 8192
rect 12256 8128 12264 8192
rect 11944 8058 11986 8128
rect 12222 8058 12264 8128
rect 11944 7104 12264 8058
rect 11944 7040 11952 7104
rect 12016 7040 12032 7104
rect 12096 7040 12112 7104
rect 12176 7040 12192 7104
rect 12256 7040 12264 7104
rect 11944 6016 12264 7040
rect 11944 5952 11952 6016
rect 12016 5952 12032 6016
rect 12096 5952 12112 6016
rect 12176 5952 12192 6016
rect 12256 5952 12264 6016
rect 11944 4928 12264 5952
rect 11944 4864 11952 4928
rect 12016 4864 12032 4928
rect 12096 4864 12112 4928
rect 12176 4864 12192 4928
rect 12256 4864 12264 4928
rect 11944 3840 12264 4864
rect 11944 3776 11952 3840
rect 12016 3776 12032 3840
rect 12096 3776 12112 3840
rect 12176 3776 12192 3840
rect 12256 3776 12264 3840
rect 11944 3294 12264 3776
rect 11944 3058 11986 3294
rect 12222 3058 12264 3294
rect 11944 2752 12264 3058
rect 11944 2688 11952 2752
rect 12016 2688 12032 2752
rect 12096 2688 12112 2752
rect 12176 2688 12192 2752
rect 12256 2688 12264 2752
rect 11944 2128 12264 2688
rect 12604 37024 12924 37584
rect 12604 36960 12612 37024
rect 12676 36960 12692 37024
rect 12756 36960 12772 37024
rect 12836 36960 12852 37024
rect 12916 36960 12924 37024
rect 12604 35936 12924 36960
rect 12604 35872 12612 35936
rect 12676 35872 12692 35936
rect 12756 35872 12772 35936
rect 12836 35872 12852 35936
rect 12916 35872 12924 35936
rect 12604 34848 12924 35872
rect 12604 34784 12612 34848
rect 12676 34784 12692 34848
rect 12756 34784 12772 34848
rect 12836 34784 12852 34848
rect 12916 34784 12924 34848
rect 12604 33954 12924 34784
rect 12604 33760 12646 33954
rect 12882 33760 12924 33954
rect 12604 33696 12612 33760
rect 12676 33696 12692 33718
rect 12756 33696 12772 33718
rect 12836 33696 12852 33718
rect 12916 33696 12924 33760
rect 12604 32672 12924 33696
rect 12604 32608 12612 32672
rect 12676 32608 12692 32672
rect 12756 32608 12772 32672
rect 12836 32608 12852 32672
rect 12916 32608 12924 32672
rect 12604 31584 12924 32608
rect 12604 31520 12612 31584
rect 12676 31520 12692 31584
rect 12756 31520 12772 31584
rect 12836 31520 12852 31584
rect 12916 31520 12924 31584
rect 12604 30496 12924 31520
rect 12604 30432 12612 30496
rect 12676 30432 12692 30496
rect 12756 30432 12772 30496
rect 12836 30432 12852 30496
rect 12916 30432 12924 30496
rect 12604 29408 12924 30432
rect 12604 29344 12612 29408
rect 12676 29344 12692 29408
rect 12756 29344 12772 29408
rect 12836 29344 12852 29408
rect 12916 29344 12924 29408
rect 12604 28954 12924 29344
rect 12604 28718 12646 28954
rect 12882 28718 12924 28954
rect 12604 28320 12924 28718
rect 12604 28256 12612 28320
rect 12676 28256 12692 28320
rect 12756 28256 12772 28320
rect 12836 28256 12852 28320
rect 12916 28256 12924 28320
rect 12604 27232 12924 28256
rect 12604 27168 12612 27232
rect 12676 27168 12692 27232
rect 12756 27168 12772 27232
rect 12836 27168 12852 27232
rect 12916 27168 12924 27232
rect 12604 26144 12924 27168
rect 12604 26080 12612 26144
rect 12676 26080 12692 26144
rect 12756 26080 12772 26144
rect 12836 26080 12852 26144
rect 12916 26080 12924 26144
rect 12604 25056 12924 26080
rect 12604 24992 12612 25056
rect 12676 24992 12692 25056
rect 12756 24992 12772 25056
rect 12836 24992 12852 25056
rect 12916 24992 12924 25056
rect 12604 23968 12924 24992
rect 12604 23904 12612 23968
rect 12676 23954 12692 23968
rect 12756 23954 12772 23968
rect 12836 23954 12852 23968
rect 12916 23904 12924 23968
rect 12604 23718 12646 23904
rect 12882 23718 12924 23904
rect 12604 22880 12924 23718
rect 12604 22816 12612 22880
rect 12676 22816 12692 22880
rect 12756 22816 12772 22880
rect 12836 22816 12852 22880
rect 12916 22816 12924 22880
rect 12604 21792 12924 22816
rect 12604 21728 12612 21792
rect 12676 21728 12692 21792
rect 12756 21728 12772 21792
rect 12836 21728 12852 21792
rect 12916 21728 12924 21792
rect 12604 20704 12924 21728
rect 12604 20640 12612 20704
rect 12676 20640 12692 20704
rect 12756 20640 12772 20704
rect 12836 20640 12852 20704
rect 12916 20640 12924 20704
rect 12604 19616 12924 20640
rect 12604 19552 12612 19616
rect 12676 19552 12692 19616
rect 12756 19552 12772 19616
rect 12836 19552 12852 19616
rect 12916 19552 12924 19616
rect 12604 18954 12924 19552
rect 12604 18718 12646 18954
rect 12882 18718 12924 18954
rect 12604 18528 12924 18718
rect 12604 18464 12612 18528
rect 12676 18464 12692 18528
rect 12756 18464 12772 18528
rect 12836 18464 12852 18528
rect 12916 18464 12924 18528
rect 12604 17440 12924 18464
rect 12604 17376 12612 17440
rect 12676 17376 12692 17440
rect 12756 17376 12772 17440
rect 12836 17376 12852 17440
rect 12916 17376 12924 17440
rect 12604 16352 12924 17376
rect 12604 16288 12612 16352
rect 12676 16288 12692 16352
rect 12756 16288 12772 16352
rect 12836 16288 12852 16352
rect 12916 16288 12924 16352
rect 12604 15264 12924 16288
rect 12604 15200 12612 15264
rect 12676 15200 12692 15264
rect 12756 15200 12772 15264
rect 12836 15200 12852 15264
rect 12916 15200 12924 15264
rect 12604 14176 12924 15200
rect 12604 14112 12612 14176
rect 12676 14112 12692 14176
rect 12756 14112 12772 14176
rect 12836 14112 12852 14176
rect 12916 14112 12924 14176
rect 12604 13954 12924 14112
rect 12604 13718 12646 13954
rect 12882 13718 12924 13954
rect 12604 13088 12924 13718
rect 12604 13024 12612 13088
rect 12676 13024 12692 13088
rect 12756 13024 12772 13088
rect 12836 13024 12852 13088
rect 12916 13024 12924 13088
rect 12604 12000 12924 13024
rect 12604 11936 12612 12000
rect 12676 11936 12692 12000
rect 12756 11936 12772 12000
rect 12836 11936 12852 12000
rect 12916 11936 12924 12000
rect 12604 10912 12924 11936
rect 12604 10848 12612 10912
rect 12676 10848 12692 10912
rect 12756 10848 12772 10912
rect 12836 10848 12852 10912
rect 12916 10848 12924 10912
rect 12604 9824 12924 10848
rect 12604 9760 12612 9824
rect 12676 9760 12692 9824
rect 12756 9760 12772 9824
rect 12836 9760 12852 9824
rect 12916 9760 12924 9824
rect 12604 8954 12924 9760
rect 12604 8736 12646 8954
rect 12882 8736 12924 8954
rect 12604 8672 12612 8736
rect 12676 8672 12692 8718
rect 12756 8672 12772 8718
rect 12836 8672 12852 8718
rect 12916 8672 12924 8736
rect 12604 7648 12924 8672
rect 12604 7584 12612 7648
rect 12676 7584 12692 7648
rect 12756 7584 12772 7648
rect 12836 7584 12852 7648
rect 12916 7584 12924 7648
rect 12604 6560 12924 7584
rect 12604 6496 12612 6560
rect 12676 6496 12692 6560
rect 12756 6496 12772 6560
rect 12836 6496 12852 6560
rect 12916 6496 12924 6560
rect 12604 5472 12924 6496
rect 12604 5408 12612 5472
rect 12676 5408 12692 5472
rect 12756 5408 12772 5472
rect 12836 5408 12852 5472
rect 12916 5408 12924 5472
rect 12604 4384 12924 5408
rect 12604 4320 12612 4384
rect 12676 4320 12692 4384
rect 12756 4320 12772 4384
rect 12836 4320 12852 4384
rect 12916 4320 12924 4384
rect 12604 3954 12924 4320
rect 12604 3718 12646 3954
rect 12882 3718 12924 3954
rect 12604 3296 12924 3718
rect 12604 3232 12612 3296
rect 12676 3232 12692 3296
rect 12756 3232 12772 3296
rect 12836 3232 12852 3296
rect 12916 3232 12924 3296
rect 12604 2208 12924 3232
rect 12604 2144 12612 2208
rect 12676 2144 12692 2208
rect 12756 2144 12772 2208
rect 12836 2144 12852 2208
rect 12916 2144 12924 2208
rect 12604 2128 12924 2144
rect 16944 37568 17264 37584
rect 16944 37504 16952 37568
rect 17016 37504 17032 37568
rect 17096 37504 17112 37568
rect 17176 37504 17192 37568
rect 17256 37504 17264 37568
rect 16944 36480 17264 37504
rect 16944 36416 16952 36480
rect 17016 36416 17032 36480
rect 17096 36416 17112 36480
rect 17176 36416 17192 36480
rect 17256 36416 17264 36480
rect 16944 35392 17264 36416
rect 16944 35328 16952 35392
rect 17016 35328 17032 35392
rect 17096 35328 17112 35392
rect 17176 35328 17192 35392
rect 17256 35328 17264 35392
rect 16944 34304 17264 35328
rect 16944 34240 16952 34304
rect 17016 34240 17032 34304
rect 17096 34240 17112 34304
rect 17176 34240 17192 34304
rect 17256 34240 17264 34304
rect 16944 33294 17264 34240
rect 16944 33216 16986 33294
rect 17222 33216 17264 33294
rect 16944 33152 16952 33216
rect 17256 33152 17264 33216
rect 16944 33058 16986 33152
rect 17222 33058 17264 33152
rect 16944 32128 17264 33058
rect 16944 32064 16952 32128
rect 17016 32064 17032 32128
rect 17096 32064 17112 32128
rect 17176 32064 17192 32128
rect 17256 32064 17264 32128
rect 16944 31040 17264 32064
rect 16944 30976 16952 31040
rect 17016 30976 17032 31040
rect 17096 30976 17112 31040
rect 17176 30976 17192 31040
rect 17256 30976 17264 31040
rect 16944 29952 17264 30976
rect 16944 29888 16952 29952
rect 17016 29888 17032 29952
rect 17096 29888 17112 29952
rect 17176 29888 17192 29952
rect 17256 29888 17264 29952
rect 16944 28864 17264 29888
rect 16944 28800 16952 28864
rect 17016 28800 17032 28864
rect 17096 28800 17112 28864
rect 17176 28800 17192 28864
rect 17256 28800 17264 28864
rect 16944 28294 17264 28800
rect 16944 28058 16986 28294
rect 17222 28058 17264 28294
rect 16944 27776 17264 28058
rect 16944 27712 16952 27776
rect 17016 27712 17032 27776
rect 17096 27712 17112 27776
rect 17176 27712 17192 27776
rect 17256 27712 17264 27776
rect 16944 26688 17264 27712
rect 16944 26624 16952 26688
rect 17016 26624 17032 26688
rect 17096 26624 17112 26688
rect 17176 26624 17192 26688
rect 17256 26624 17264 26688
rect 16944 25600 17264 26624
rect 16944 25536 16952 25600
rect 17016 25536 17032 25600
rect 17096 25536 17112 25600
rect 17176 25536 17192 25600
rect 17256 25536 17264 25600
rect 16944 24512 17264 25536
rect 16944 24448 16952 24512
rect 17016 24448 17032 24512
rect 17096 24448 17112 24512
rect 17176 24448 17192 24512
rect 17256 24448 17264 24512
rect 16944 23424 17264 24448
rect 16944 23360 16952 23424
rect 17016 23360 17032 23424
rect 17096 23360 17112 23424
rect 17176 23360 17192 23424
rect 17256 23360 17264 23424
rect 16944 23294 17264 23360
rect 16944 23058 16986 23294
rect 17222 23058 17264 23294
rect 16944 22336 17264 23058
rect 16944 22272 16952 22336
rect 17016 22272 17032 22336
rect 17096 22272 17112 22336
rect 17176 22272 17192 22336
rect 17256 22272 17264 22336
rect 16944 21248 17264 22272
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 18294 17264 19008
rect 16944 18058 16986 18294
rect 17222 18058 17264 18294
rect 16944 17984 17264 18058
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13294 17264 13568
rect 16944 13058 16986 13294
rect 17222 13058 17264 13294
rect 16944 12544 17264 13058
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8294 17264 9216
rect 16944 8192 16986 8294
rect 17222 8192 17264 8294
rect 16944 8128 16952 8192
rect 17256 8128 17264 8192
rect 16944 8058 16986 8128
rect 17222 8058 17264 8128
rect 16944 7104 17264 8058
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3294 17264 3776
rect 16944 3058 16986 3294
rect 17222 3058 17264 3294
rect 16944 2752 17264 3058
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 17604 37024 17924 37584
rect 17604 36960 17612 37024
rect 17676 36960 17692 37024
rect 17756 36960 17772 37024
rect 17836 36960 17852 37024
rect 17916 36960 17924 37024
rect 17604 35936 17924 36960
rect 17604 35872 17612 35936
rect 17676 35872 17692 35936
rect 17756 35872 17772 35936
rect 17836 35872 17852 35936
rect 17916 35872 17924 35936
rect 17604 34848 17924 35872
rect 17604 34784 17612 34848
rect 17676 34784 17692 34848
rect 17756 34784 17772 34848
rect 17836 34784 17852 34848
rect 17916 34784 17924 34848
rect 17604 33954 17924 34784
rect 17604 33760 17646 33954
rect 17882 33760 17924 33954
rect 17604 33696 17612 33760
rect 17676 33696 17692 33718
rect 17756 33696 17772 33718
rect 17836 33696 17852 33718
rect 17916 33696 17924 33760
rect 17604 32672 17924 33696
rect 17604 32608 17612 32672
rect 17676 32608 17692 32672
rect 17756 32608 17772 32672
rect 17836 32608 17852 32672
rect 17916 32608 17924 32672
rect 17604 31584 17924 32608
rect 17604 31520 17612 31584
rect 17676 31520 17692 31584
rect 17756 31520 17772 31584
rect 17836 31520 17852 31584
rect 17916 31520 17924 31584
rect 17604 30496 17924 31520
rect 17604 30432 17612 30496
rect 17676 30432 17692 30496
rect 17756 30432 17772 30496
rect 17836 30432 17852 30496
rect 17916 30432 17924 30496
rect 17604 29408 17924 30432
rect 17604 29344 17612 29408
rect 17676 29344 17692 29408
rect 17756 29344 17772 29408
rect 17836 29344 17852 29408
rect 17916 29344 17924 29408
rect 17604 28954 17924 29344
rect 17604 28718 17646 28954
rect 17882 28718 17924 28954
rect 17604 28320 17924 28718
rect 17604 28256 17612 28320
rect 17676 28256 17692 28320
rect 17756 28256 17772 28320
rect 17836 28256 17852 28320
rect 17916 28256 17924 28320
rect 17604 27232 17924 28256
rect 17604 27168 17612 27232
rect 17676 27168 17692 27232
rect 17756 27168 17772 27232
rect 17836 27168 17852 27232
rect 17916 27168 17924 27232
rect 17604 26144 17924 27168
rect 17604 26080 17612 26144
rect 17676 26080 17692 26144
rect 17756 26080 17772 26144
rect 17836 26080 17852 26144
rect 17916 26080 17924 26144
rect 17604 25056 17924 26080
rect 17604 24992 17612 25056
rect 17676 24992 17692 25056
rect 17756 24992 17772 25056
rect 17836 24992 17852 25056
rect 17916 24992 17924 25056
rect 17604 23968 17924 24992
rect 17604 23904 17612 23968
rect 17676 23954 17692 23968
rect 17756 23954 17772 23968
rect 17836 23954 17852 23968
rect 17916 23904 17924 23968
rect 17604 23718 17646 23904
rect 17882 23718 17924 23904
rect 17604 22880 17924 23718
rect 17604 22816 17612 22880
rect 17676 22816 17692 22880
rect 17756 22816 17772 22880
rect 17836 22816 17852 22880
rect 17916 22816 17924 22880
rect 17604 21792 17924 22816
rect 17604 21728 17612 21792
rect 17676 21728 17692 21792
rect 17756 21728 17772 21792
rect 17836 21728 17852 21792
rect 17916 21728 17924 21792
rect 17604 20704 17924 21728
rect 17604 20640 17612 20704
rect 17676 20640 17692 20704
rect 17756 20640 17772 20704
rect 17836 20640 17852 20704
rect 17916 20640 17924 20704
rect 17604 19616 17924 20640
rect 17604 19552 17612 19616
rect 17676 19552 17692 19616
rect 17756 19552 17772 19616
rect 17836 19552 17852 19616
rect 17916 19552 17924 19616
rect 17604 18954 17924 19552
rect 17604 18718 17646 18954
rect 17882 18718 17924 18954
rect 17604 18528 17924 18718
rect 17604 18464 17612 18528
rect 17676 18464 17692 18528
rect 17756 18464 17772 18528
rect 17836 18464 17852 18528
rect 17916 18464 17924 18528
rect 17604 17440 17924 18464
rect 17604 17376 17612 17440
rect 17676 17376 17692 17440
rect 17756 17376 17772 17440
rect 17836 17376 17852 17440
rect 17916 17376 17924 17440
rect 17604 16352 17924 17376
rect 17604 16288 17612 16352
rect 17676 16288 17692 16352
rect 17756 16288 17772 16352
rect 17836 16288 17852 16352
rect 17916 16288 17924 16352
rect 17604 15264 17924 16288
rect 17604 15200 17612 15264
rect 17676 15200 17692 15264
rect 17756 15200 17772 15264
rect 17836 15200 17852 15264
rect 17916 15200 17924 15264
rect 17604 14176 17924 15200
rect 17604 14112 17612 14176
rect 17676 14112 17692 14176
rect 17756 14112 17772 14176
rect 17836 14112 17852 14176
rect 17916 14112 17924 14176
rect 17604 13954 17924 14112
rect 17604 13718 17646 13954
rect 17882 13718 17924 13954
rect 17604 13088 17924 13718
rect 17604 13024 17612 13088
rect 17676 13024 17692 13088
rect 17756 13024 17772 13088
rect 17836 13024 17852 13088
rect 17916 13024 17924 13088
rect 17604 12000 17924 13024
rect 17604 11936 17612 12000
rect 17676 11936 17692 12000
rect 17756 11936 17772 12000
rect 17836 11936 17852 12000
rect 17916 11936 17924 12000
rect 17604 10912 17924 11936
rect 17604 10848 17612 10912
rect 17676 10848 17692 10912
rect 17756 10848 17772 10912
rect 17836 10848 17852 10912
rect 17916 10848 17924 10912
rect 17604 9824 17924 10848
rect 17604 9760 17612 9824
rect 17676 9760 17692 9824
rect 17756 9760 17772 9824
rect 17836 9760 17852 9824
rect 17916 9760 17924 9824
rect 17604 8954 17924 9760
rect 17604 8736 17646 8954
rect 17882 8736 17924 8954
rect 17604 8672 17612 8736
rect 17676 8672 17692 8718
rect 17756 8672 17772 8718
rect 17836 8672 17852 8718
rect 17916 8672 17924 8736
rect 17604 7648 17924 8672
rect 17604 7584 17612 7648
rect 17676 7584 17692 7648
rect 17756 7584 17772 7648
rect 17836 7584 17852 7648
rect 17916 7584 17924 7648
rect 17604 6560 17924 7584
rect 17604 6496 17612 6560
rect 17676 6496 17692 6560
rect 17756 6496 17772 6560
rect 17836 6496 17852 6560
rect 17916 6496 17924 6560
rect 17604 5472 17924 6496
rect 17604 5408 17612 5472
rect 17676 5408 17692 5472
rect 17756 5408 17772 5472
rect 17836 5408 17852 5472
rect 17916 5408 17924 5472
rect 17604 4384 17924 5408
rect 17604 4320 17612 4384
rect 17676 4320 17692 4384
rect 17756 4320 17772 4384
rect 17836 4320 17852 4384
rect 17916 4320 17924 4384
rect 17604 3954 17924 4320
rect 17604 3718 17646 3954
rect 17882 3718 17924 3954
rect 17604 3296 17924 3718
rect 17604 3232 17612 3296
rect 17676 3232 17692 3296
rect 17756 3232 17772 3296
rect 17836 3232 17852 3296
rect 17916 3232 17924 3296
rect 17604 2208 17924 3232
rect 17604 2144 17612 2208
rect 17676 2144 17692 2208
rect 17756 2144 17772 2208
rect 17836 2144 17852 2208
rect 17916 2144 17924 2208
rect 17604 2128 17924 2144
rect 21944 37568 22264 37584
rect 21944 37504 21952 37568
rect 22016 37504 22032 37568
rect 22096 37504 22112 37568
rect 22176 37504 22192 37568
rect 22256 37504 22264 37568
rect 21944 36480 22264 37504
rect 21944 36416 21952 36480
rect 22016 36416 22032 36480
rect 22096 36416 22112 36480
rect 22176 36416 22192 36480
rect 22256 36416 22264 36480
rect 21944 35392 22264 36416
rect 21944 35328 21952 35392
rect 22016 35328 22032 35392
rect 22096 35328 22112 35392
rect 22176 35328 22192 35392
rect 22256 35328 22264 35392
rect 21944 34304 22264 35328
rect 21944 34240 21952 34304
rect 22016 34240 22032 34304
rect 22096 34240 22112 34304
rect 22176 34240 22192 34304
rect 22256 34240 22264 34304
rect 21944 33294 22264 34240
rect 21944 33216 21986 33294
rect 22222 33216 22264 33294
rect 21944 33152 21952 33216
rect 22256 33152 22264 33216
rect 21944 33058 21986 33152
rect 22222 33058 22264 33152
rect 21944 32128 22264 33058
rect 21944 32064 21952 32128
rect 22016 32064 22032 32128
rect 22096 32064 22112 32128
rect 22176 32064 22192 32128
rect 22256 32064 22264 32128
rect 21944 31040 22264 32064
rect 21944 30976 21952 31040
rect 22016 30976 22032 31040
rect 22096 30976 22112 31040
rect 22176 30976 22192 31040
rect 22256 30976 22264 31040
rect 21944 29952 22264 30976
rect 21944 29888 21952 29952
rect 22016 29888 22032 29952
rect 22096 29888 22112 29952
rect 22176 29888 22192 29952
rect 22256 29888 22264 29952
rect 21944 28864 22264 29888
rect 21944 28800 21952 28864
rect 22016 28800 22032 28864
rect 22096 28800 22112 28864
rect 22176 28800 22192 28864
rect 22256 28800 22264 28864
rect 21944 28294 22264 28800
rect 21944 28058 21986 28294
rect 22222 28058 22264 28294
rect 21944 27776 22264 28058
rect 21944 27712 21952 27776
rect 22016 27712 22032 27776
rect 22096 27712 22112 27776
rect 22176 27712 22192 27776
rect 22256 27712 22264 27776
rect 21944 26688 22264 27712
rect 21944 26624 21952 26688
rect 22016 26624 22032 26688
rect 22096 26624 22112 26688
rect 22176 26624 22192 26688
rect 22256 26624 22264 26688
rect 21944 25600 22264 26624
rect 21944 25536 21952 25600
rect 22016 25536 22032 25600
rect 22096 25536 22112 25600
rect 22176 25536 22192 25600
rect 22256 25536 22264 25600
rect 21944 24512 22264 25536
rect 21944 24448 21952 24512
rect 22016 24448 22032 24512
rect 22096 24448 22112 24512
rect 22176 24448 22192 24512
rect 22256 24448 22264 24512
rect 21944 23424 22264 24448
rect 21944 23360 21952 23424
rect 22016 23360 22032 23424
rect 22096 23360 22112 23424
rect 22176 23360 22192 23424
rect 22256 23360 22264 23424
rect 21944 23294 22264 23360
rect 21944 23058 21986 23294
rect 22222 23058 22264 23294
rect 21944 22336 22264 23058
rect 21944 22272 21952 22336
rect 22016 22272 22032 22336
rect 22096 22272 22112 22336
rect 22176 22272 22192 22336
rect 22256 22272 22264 22336
rect 21944 21248 22264 22272
rect 21944 21184 21952 21248
rect 22016 21184 22032 21248
rect 22096 21184 22112 21248
rect 22176 21184 22192 21248
rect 22256 21184 22264 21248
rect 21944 20160 22264 21184
rect 21944 20096 21952 20160
rect 22016 20096 22032 20160
rect 22096 20096 22112 20160
rect 22176 20096 22192 20160
rect 22256 20096 22264 20160
rect 21944 19072 22264 20096
rect 21944 19008 21952 19072
rect 22016 19008 22032 19072
rect 22096 19008 22112 19072
rect 22176 19008 22192 19072
rect 22256 19008 22264 19072
rect 21944 18294 22264 19008
rect 21944 18058 21986 18294
rect 22222 18058 22264 18294
rect 21944 17984 22264 18058
rect 21944 17920 21952 17984
rect 22016 17920 22032 17984
rect 22096 17920 22112 17984
rect 22176 17920 22192 17984
rect 22256 17920 22264 17984
rect 21944 16896 22264 17920
rect 21944 16832 21952 16896
rect 22016 16832 22032 16896
rect 22096 16832 22112 16896
rect 22176 16832 22192 16896
rect 22256 16832 22264 16896
rect 21944 15808 22264 16832
rect 21944 15744 21952 15808
rect 22016 15744 22032 15808
rect 22096 15744 22112 15808
rect 22176 15744 22192 15808
rect 22256 15744 22264 15808
rect 21944 14720 22264 15744
rect 21944 14656 21952 14720
rect 22016 14656 22032 14720
rect 22096 14656 22112 14720
rect 22176 14656 22192 14720
rect 22256 14656 22264 14720
rect 21944 13632 22264 14656
rect 21944 13568 21952 13632
rect 22016 13568 22032 13632
rect 22096 13568 22112 13632
rect 22176 13568 22192 13632
rect 22256 13568 22264 13632
rect 21944 13294 22264 13568
rect 21944 13058 21986 13294
rect 22222 13058 22264 13294
rect 21944 12544 22264 13058
rect 21944 12480 21952 12544
rect 22016 12480 22032 12544
rect 22096 12480 22112 12544
rect 22176 12480 22192 12544
rect 22256 12480 22264 12544
rect 21944 11456 22264 12480
rect 21944 11392 21952 11456
rect 22016 11392 22032 11456
rect 22096 11392 22112 11456
rect 22176 11392 22192 11456
rect 22256 11392 22264 11456
rect 21944 10368 22264 11392
rect 21944 10304 21952 10368
rect 22016 10304 22032 10368
rect 22096 10304 22112 10368
rect 22176 10304 22192 10368
rect 22256 10304 22264 10368
rect 21944 9280 22264 10304
rect 21944 9216 21952 9280
rect 22016 9216 22032 9280
rect 22096 9216 22112 9280
rect 22176 9216 22192 9280
rect 22256 9216 22264 9280
rect 21944 8294 22264 9216
rect 21944 8192 21986 8294
rect 22222 8192 22264 8294
rect 21944 8128 21952 8192
rect 22256 8128 22264 8192
rect 21944 8058 21986 8128
rect 22222 8058 22264 8128
rect 21944 7104 22264 8058
rect 21944 7040 21952 7104
rect 22016 7040 22032 7104
rect 22096 7040 22112 7104
rect 22176 7040 22192 7104
rect 22256 7040 22264 7104
rect 21944 6016 22264 7040
rect 21944 5952 21952 6016
rect 22016 5952 22032 6016
rect 22096 5952 22112 6016
rect 22176 5952 22192 6016
rect 22256 5952 22264 6016
rect 21944 4928 22264 5952
rect 21944 4864 21952 4928
rect 22016 4864 22032 4928
rect 22096 4864 22112 4928
rect 22176 4864 22192 4928
rect 22256 4864 22264 4928
rect 21944 3840 22264 4864
rect 21944 3776 21952 3840
rect 22016 3776 22032 3840
rect 22096 3776 22112 3840
rect 22176 3776 22192 3840
rect 22256 3776 22264 3840
rect 21944 3294 22264 3776
rect 21944 3058 21986 3294
rect 22222 3058 22264 3294
rect 21944 2752 22264 3058
rect 21944 2688 21952 2752
rect 22016 2688 22032 2752
rect 22096 2688 22112 2752
rect 22176 2688 22192 2752
rect 22256 2688 22264 2752
rect 21944 2128 22264 2688
rect 22604 37024 22924 37584
rect 22604 36960 22612 37024
rect 22676 36960 22692 37024
rect 22756 36960 22772 37024
rect 22836 36960 22852 37024
rect 22916 36960 22924 37024
rect 22604 35936 22924 36960
rect 22604 35872 22612 35936
rect 22676 35872 22692 35936
rect 22756 35872 22772 35936
rect 22836 35872 22852 35936
rect 22916 35872 22924 35936
rect 22604 34848 22924 35872
rect 22604 34784 22612 34848
rect 22676 34784 22692 34848
rect 22756 34784 22772 34848
rect 22836 34784 22852 34848
rect 22916 34784 22924 34848
rect 22604 33954 22924 34784
rect 22604 33760 22646 33954
rect 22882 33760 22924 33954
rect 22604 33696 22612 33760
rect 22676 33696 22692 33718
rect 22756 33696 22772 33718
rect 22836 33696 22852 33718
rect 22916 33696 22924 33760
rect 22604 32672 22924 33696
rect 22604 32608 22612 32672
rect 22676 32608 22692 32672
rect 22756 32608 22772 32672
rect 22836 32608 22852 32672
rect 22916 32608 22924 32672
rect 22604 31584 22924 32608
rect 22604 31520 22612 31584
rect 22676 31520 22692 31584
rect 22756 31520 22772 31584
rect 22836 31520 22852 31584
rect 22916 31520 22924 31584
rect 22604 30496 22924 31520
rect 22604 30432 22612 30496
rect 22676 30432 22692 30496
rect 22756 30432 22772 30496
rect 22836 30432 22852 30496
rect 22916 30432 22924 30496
rect 22604 29408 22924 30432
rect 22604 29344 22612 29408
rect 22676 29344 22692 29408
rect 22756 29344 22772 29408
rect 22836 29344 22852 29408
rect 22916 29344 22924 29408
rect 22604 28954 22924 29344
rect 22604 28718 22646 28954
rect 22882 28718 22924 28954
rect 22604 28320 22924 28718
rect 22604 28256 22612 28320
rect 22676 28256 22692 28320
rect 22756 28256 22772 28320
rect 22836 28256 22852 28320
rect 22916 28256 22924 28320
rect 22604 27232 22924 28256
rect 22604 27168 22612 27232
rect 22676 27168 22692 27232
rect 22756 27168 22772 27232
rect 22836 27168 22852 27232
rect 22916 27168 22924 27232
rect 22604 26144 22924 27168
rect 22604 26080 22612 26144
rect 22676 26080 22692 26144
rect 22756 26080 22772 26144
rect 22836 26080 22852 26144
rect 22916 26080 22924 26144
rect 22604 25056 22924 26080
rect 22604 24992 22612 25056
rect 22676 24992 22692 25056
rect 22756 24992 22772 25056
rect 22836 24992 22852 25056
rect 22916 24992 22924 25056
rect 22604 23968 22924 24992
rect 22604 23904 22612 23968
rect 22676 23954 22692 23968
rect 22756 23954 22772 23968
rect 22836 23954 22852 23968
rect 22916 23904 22924 23968
rect 22604 23718 22646 23904
rect 22882 23718 22924 23904
rect 22604 22880 22924 23718
rect 22604 22816 22612 22880
rect 22676 22816 22692 22880
rect 22756 22816 22772 22880
rect 22836 22816 22852 22880
rect 22916 22816 22924 22880
rect 22604 21792 22924 22816
rect 22604 21728 22612 21792
rect 22676 21728 22692 21792
rect 22756 21728 22772 21792
rect 22836 21728 22852 21792
rect 22916 21728 22924 21792
rect 22604 20704 22924 21728
rect 22604 20640 22612 20704
rect 22676 20640 22692 20704
rect 22756 20640 22772 20704
rect 22836 20640 22852 20704
rect 22916 20640 22924 20704
rect 22604 19616 22924 20640
rect 22604 19552 22612 19616
rect 22676 19552 22692 19616
rect 22756 19552 22772 19616
rect 22836 19552 22852 19616
rect 22916 19552 22924 19616
rect 22604 18954 22924 19552
rect 22604 18718 22646 18954
rect 22882 18718 22924 18954
rect 22604 18528 22924 18718
rect 22604 18464 22612 18528
rect 22676 18464 22692 18528
rect 22756 18464 22772 18528
rect 22836 18464 22852 18528
rect 22916 18464 22924 18528
rect 22604 17440 22924 18464
rect 22604 17376 22612 17440
rect 22676 17376 22692 17440
rect 22756 17376 22772 17440
rect 22836 17376 22852 17440
rect 22916 17376 22924 17440
rect 22604 16352 22924 17376
rect 22604 16288 22612 16352
rect 22676 16288 22692 16352
rect 22756 16288 22772 16352
rect 22836 16288 22852 16352
rect 22916 16288 22924 16352
rect 22604 15264 22924 16288
rect 22604 15200 22612 15264
rect 22676 15200 22692 15264
rect 22756 15200 22772 15264
rect 22836 15200 22852 15264
rect 22916 15200 22924 15264
rect 22604 14176 22924 15200
rect 22604 14112 22612 14176
rect 22676 14112 22692 14176
rect 22756 14112 22772 14176
rect 22836 14112 22852 14176
rect 22916 14112 22924 14176
rect 22604 13954 22924 14112
rect 22604 13718 22646 13954
rect 22882 13718 22924 13954
rect 22604 13088 22924 13718
rect 22604 13024 22612 13088
rect 22676 13024 22692 13088
rect 22756 13024 22772 13088
rect 22836 13024 22852 13088
rect 22916 13024 22924 13088
rect 22604 12000 22924 13024
rect 22604 11936 22612 12000
rect 22676 11936 22692 12000
rect 22756 11936 22772 12000
rect 22836 11936 22852 12000
rect 22916 11936 22924 12000
rect 22604 10912 22924 11936
rect 22604 10848 22612 10912
rect 22676 10848 22692 10912
rect 22756 10848 22772 10912
rect 22836 10848 22852 10912
rect 22916 10848 22924 10912
rect 22604 9824 22924 10848
rect 22604 9760 22612 9824
rect 22676 9760 22692 9824
rect 22756 9760 22772 9824
rect 22836 9760 22852 9824
rect 22916 9760 22924 9824
rect 22604 8954 22924 9760
rect 22604 8736 22646 8954
rect 22882 8736 22924 8954
rect 22604 8672 22612 8736
rect 22676 8672 22692 8718
rect 22756 8672 22772 8718
rect 22836 8672 22852 8718
rect 22916 8672 22924 8736
rect 22604 7648 22924 8672
rect 22604 7584 22612 7648
rect 22676 7584 22692 7648
rect 22756 7584 22772 7648
rect 22836 7584 22852 7648
rect 22916 7584 22924 7648
rect 22604 6560 22924 7584
rect 22604 6496 22612 6560
rect 22676 6496 22692 6560
rect 22756 6496 22772 6560
rect 22836 6496 22852 6560
rect 22916 6496 22924 6560
rect 22604 5472 22924 6496
rect 22604 5408 22612 5472
rect 22676 5408 22692 5472
rect 22756 5408 22772 5472
rect 22836 5408 22852 5472
rect 22916 5408 22924 5472
rect 22604 4384 22924 5408
rect 22604 4320 22612 4384
rect 22676 4320 22692 4384
rect 22756 4320 22772 4384
rect 22836 4320 22852 4384
rect 22916 4320 22924 4384
rect 22604 3954 22924 4320
rect 22604 3718 22646 3954
rect 22882 3718 22924 3954
rect 22604 3296 22924 3718
rect 22604 3232 22612 3296
rect 22676 3232 22692 3296
rect 22756 3232 22772 3296
rect 22836 3232 22852 3296
rect 22916 3232 22924 3296
rect 22604 2208 22924 3232
rect 22604 2144 22612 2208
rect 22676 2144 22692 2208
rect 22756 2144 22772 2208
rect 22836 2144 22852 2208
rect 22916 2144 22924 2208
rect 22604 2128 22924 2144
rect 26944 37568 27264 37584
rect 26944 37504 26952 37568
rect 27016 37504 27032 37568
rect 27096 37504 27112 37568
rect 27176 37504 27192 37568
rect 27256 37504 27264 37568
rect 26944 36480 27264 37504
rect 26944 36416 26952 36480
rect 27016 36416 27032 36480
rect 27096 36416 27112 36480
rect 27176 36416 27192 36480
rect 27256 36416 27264 36480
rect 26944 35392 27264 36416
rect 26944 35328 26952 35392
rect 27016 35328 27032 35392
rect 27096 35328 27112 35392
rect 27176 35328 27192 35392
rect 27256 35328 27264 35392
rect 26944 34304 27264 35328
rect 26944 34240 26952 34304
rect 27016 34240 27032 34304
rect 27096 34240 27112 34304
rect 27176 34240 27192 34304
rect 27256 34240 27264 34304
rect 26944 33294 27264 34240
rect 26944 33216 26986 33294
rect 27222 33216 27264 33294
rect 26944 33152 26952 33216
rect 27256 33152 27264 33216
rect 26944 33058 26986 33152
rect 27222 33058 27264 33152
rect 26944 32128 27264 33058
rect 26944 32064 26952 32128
rect 27016 32064 27032 32128
rect 27096 32064 27112 32128
rect 27176 32064 27192 32128
rect 27256 32064 27264 32128
rect 26944 31040 27264 32064
rect 26944 30976 26952 31040
rect 27016 30976 27032 31040
rect 27096 30976 27112 31040
rect 27176 30976 27192 31040
rect 27256 30976 27264 31040
rect 26944 29952 27264 30976
rect 26944 29888 26952 29952
rect 27016 29888 27032 29952
rect 27096 29888 27112 29952
rect 27176 29888 27192 29952
rect 27256 29888 27264 29952
rect 26944 28864 27264 29888
rect 26944 28800 26952 28864
rect 27016 28800 27032 28864
rect 27096 28800 27112 28864
rect 27176 28800 27192 28864
rect 27256 28800 27264 28864
rect 26944 28294 27264 28800
rect 26944 28058 26986 28294
rect 27222 28058 27264 28294
rect 26944 27776 27264 28058
rect 26944 27712 26952 27776
rect 27016 27712 27032 27776
rect 27096 27712 27112 27776
rect 27176 27712 27192 27776
rect 27256 27712 27264 27776
rect 26944 26688 27264 27712
rect 26944 26624 26952 26688
rect 27016 26624 27032 26688
rect 27096 26624 27112 26688
rect 27176 26624 27192 26688
rect 27256 26624 27264 26688
rect 26944 25600 27264 26624
rect 26944 25536 26952 25600
rect 27016 25536 27032 25600
rect 27096 25536 27112 25600
rect 27176 25536 27192 25600
rect 27256 25536 27264 25600
rect 26944 24512 27264 25536
rect 26944 24448 26952 24512
rect 27016 24448 27032 24512
rect 27096 24448 27112 24512
rect 27176 24448 27192 24512
rect 27256 24448 27264 24512
rect 26944 23424 27264 24448
rect 26944 23360 26952 23424
rect 27016 23360 27032 23424
rect 27096 23360 27112 23424
rect 27176 23360 27192 23424
rect 27256 23360 27264 23424
rect 26944 23294 27264 23360
rect 26944 23058 26986 23294
rect 27222 23058 27264 23294
rect 26944 22336 27264 23058
rect 26944 22272 26952 22336
rect 27016 22272 27032 22336
rect 27096 22272 27112 22336
rect 27176 22272 27192 22336
rect 27256 22272 27264 22336
rect 26944 21248 27264 22272
rect 26944 21184 26952 21248
rect 27016 21184 27032 21248
rect 27096 21184 27112 21248
rect 27176 21184 27192 21248
rect 27256 21184 27264 21248
rect 26944 20160 27264 21184
rect 26944 20096 26952 20160
rect 27016 20096 27032 20160
rect 27096 20096 27112 20160
rect 27176 20096 27192 20160
rect 27256 20096 27264 20160
rect 26944 19072 27264 20096
rect 26944 19008 26952 19072
rect 27016 19008 27032 19072
rect 27096 19008 27112 19072
rect 27176 19008 27192 19072
rect 27256 19008 27264 19072
rect 26944 18294 27264 19008
rect 26944 18058 26986 18294
rect 27222 18058 27264 18294
rect 26944 17984 27264 18058
rect 26944 17920 26952 17984
rect 27016 17920 27032 17984
rect 27096 17920 27112 17984
rect 27176 17920 27192 17984
rect 27256 17920 27264 17984
rect 26944 16896 27264 17920
rect 26944 16832 26952 16896
rect 27016 16832 27032 16896
rect 27096 16832 27112 16896
rect 27176 16832 27192 16896
rect 27256 16832 27264 16896
rect 26944 15808 27264 16832
rect 26944 15744 26952 15808
rect 27016 15744 27032 15808
rect 27096 15744 27112 15808
rect 27176 15744 27192 15808
rect 27256 15744 27264 15808
rect 26944 14720 27264 15744
rect 26944 14656 26952 14720
rect 27016 14656 27032 14720
rect 27096 14656 27112 14720
rect 27176 14656 27192 14720
rect 27256 14656 27264 14720
rect 26944 13632 27264 14656
rect 26944 13568 26952 13632
rect 27016 13568 27032 13632
rect 27096 13568 27112 13632
rect 27176 13568 27192 13632
rect 27256 13568 27264 13632
rect 26944 13294 27264 13568
rect 26944 13058 26986 13294
rect 27222 13058 27264 13294
rect 26944 12544 27264 13058
rect 26944 12480 26952 12544
rect 27016 12480 27032 12544
rect 27096 12480 27112 12544
rect 27176 12480 27192 12544
rect 27256 12480 27264 12544
rect 26944 11456 27264 12480
rect 26944 11392 26952 11456
rect 27016 11392 27032 11456
rect 27096 11392 27112 11456
rect 27176 11392 27192 11456
rect 27256 11392 27264 11456
rect 26944 10368 27264 11392
rect 26944 10304 26952 10368
rect 27016 10304 27032 10368
rect 27096 10304 27112 10368
rect 27176 10304 27192 10368
rect 27256 10304 27264 10368
rect 26944 9280 27264 10304
rect 26944 9216 26952 9280
rect 27016 9216 27032 9280
rect 27096 9216 27112 9280
rect 27176 9216 27192 9280
rect 27256 9216 27264 9280
rect 26944 8294 27264 9216
rect 26944 8192 26986 8294
rect 27222 8192 27264 8294
rect 26944 8128 26952 8192
rect 27256 8128 27264 8192
rect 26944 8058 26986 8128
rect 27222 8058 27264 8128
rect 26944 7104 27264 8058
rect 26944 7040 26952 7104
rect 27016 7040 27032 7104
rect 27096 7040 27112 7104
rect 27176 7040 27192 7104
rect 27256 7040 27264 7104
rect 26944 6016 27264 7040
rect 26944 5952 26952 6016
rect 27016 5952 27032 6016
rect 27096 5952 27112 6016
rect 27176 5952 27192 6016
rect 27256 5952 27264 6016
rect 26944 4928 27264 5952
rect 26944 4864 26952 4928
rect 27016 4864 27032 4928
rect 27096 4864 27112 4928
rect 27176 4864 27192 4928
rect 27256 4864 27264 4928
rect 26944 3840 27264 4864
rect 26944 3776 26952 3840
rect 27016 3776 27032 3840
rect 27096 3776 27112 3840
rect 27176 3776 27192 3840
rect 27256 3776 27264 3840
rect 26944 3294 27264 3776
rect 26944 3058 26986 3294
rect 27222 3058 27264 3294
rect 26944 2752 27264 3058
rect 26944 2688 26952 2752
rect 27016 2688 27032 2752
rect 27096 2688 27112 2752
rect 27176 2688 27192 2752
rect 27256 2688 27264 2752
rect 26944 2128 27264 2688
rect 27604 37024 27924 37584
rect 27604 36960 27612 37024
rect 27676 36960 27692 37024
rect 27756 36960 27772 37024
rect 27836 36960 27852 37024
rect 27916 36960 27924 37024
rect 27604 35936 27924 36960
rect 27604 35872 27612 35936
rect 27676 35872 27692 35936
rect 27756 35872 27772 35936
rect 27836 35872 27852 35936
rect 27916 35872 27924 35936
rect 27604 34848 27924 35872
rect 27604 34784 27612 34848
rect 27676 34784 27692 34848
rect 27756 34784 27772 34848
rect 27836 34784 27852 34848
rect 27916 34784 27924 34848
rect 27604 33954 27924 34784
rect 27604 33760 27646 33954
rect 27882 33760 27924 33954
rect 27604 33696 27612 33760
rect 27676 33696 27692 33718
rect 27756 33696 27772 33718
rect 27836 33696 27852 33718
rect 27916 33696 27924 33760
rect 27604 32672 27924 33696
rect 27604 32608 27612 32672
rect 27676 32608 27692 32672
rect 27756 32608 27772 32672
rect 27836 32608 27852 32672
rect 27916 32608 27924 32672
rect 27604 31584 27924 32608
rect 27604 31520 27612 31584
rect 27676 31520 27692 31584
rect 27756 31520 27772 31584
rect 27836 31520 27852 31584
rect 27916 31520 27924 31584
rect 27604 30496 27924 31520
rect 27604 30432 27612 30496
rect 27676 30432 27692 30496
rect 27756 30432 27772 30496
rect 27836 30432 27852 30496
rect 27916 30432 27924 30496
rect 27604 29408 27924 30432
rect 27604 29344 27612 29408
rect 27676 29344 27692 29408
rect 27756 29344 27772 29408
rect 27836 29344 27852 29408
rect 27916 29344 27924 29408
rect 27604 28954 27924 29344
rect 27604 28718 27646 28954
rect 27882 28718 27924 28954
rect 27604 28320 27924 28718
rect 27604 28256 27612 28320
rect 27676 28256 27692 28320
rect 27756 28256 27772 28320
rect 27836 28256 27852 28320
rect 27916 28256 27924 28320
rect 27604 27232 27924 28256
rect 27604 27168 27612 27232
rect 27676 27168 27692 27232
rect 27756 27168 27772 27232
rect 27836 27168 27852 27232
rect 27916 27168 27924 27232
rect 27604 26144 27924 27168
rect 27604 26080 27612 26144
rect 27676 26080 27692 26144
rect 27756 26080 27772 26144
rect 27836 26080 27852 26144
rect 27916 26080 27924 26144
rect 27604 25056 27924 26080
rect 27604 24992 27612 25056
rect 27676 24992 27692 25056
rect 27756 24992 27772 25056
rect 27836 24992 27852 25056
rect 27916 24992 27924 25056
rect 27604 23968 27924 24992
rect 27604 23904 27612 23968
rect 27676 23954 27692 23968
rect 27756 23954 27772 23968
rect 27836 23954 27852 23968
rect 27916 23904 27924 23968
rect 27604 23718 27646 23904
rect 27882 23718 27924 23904
rect 27604 22880 27924 23718
rect 27604 22816 27612 22880
rect 27676 22816 27692 22880
rect 27756 22816 27772 22880
rect 27836 22816 27852 22880
rect 27916 22816 27924 22880
rect 27604 21792 27924 22816
rect 27604 21728 27612 21792
rect 27676 21728 27692 21792
rect 27756 21728 27772 21792
rect 27836 21728 27852 21792
rect 27916 21728 27924 21792
rect 27604 20704 27924 21728
rect 27604 20640 27612 20704
rect 27676 20640 27692 20704
rect 27756 20640 27772 20704
rect 27836 20640 27852 20704
rect 27916 20640 27924 20704
rect 27604 19616 27924 20640
rect 27604 19552 27612 19616
rect 27676 19552 27692 19616
rect 27756 19552 27772 19616
rect 27836 19552 27852 19616
rect 27916 19552 27924 19616
rect 27604 18954 27924 19552
rect 27604 18718 27646 18954
rect 27882 18718 27924 18954
rect 27604 18528 27924 18718
rect 27604 18464 27612 18528
rect 27676 18464 27692 18528
rect 27756 18464 27772 18528
rect 27836 18464 27852 18528
rect 27916 18464 27924 18528
rect 27604 17440 27924 18464
rect 27604 17376 27612 17440
rect 27676 17376 27692 17440
rect 27756 17376 27772 17440
rect 27836 17376 27852 17440
rect 27916 17376 27924 17440
rect 27604 16352 27924 17376
rect 27604 16288 27612 16352
rect 27676 16288 27692 16352
rect 27756 16288 27772 16352
rect 27836 16288 27852 16352
rect 27916 16288 27924 16352
rect 27604 15264 27924 16288
rect 27604 15200 27612 15264
rect 27676 15200 27692 15264
rect 27756 15200 27772 15264
rect 27836 15200 27852 15264
rect 27916 15200 27924 15264
rect 27604 14176 27924 15200
rect 27604 14112 27612 14176
rect 27676 14112 27692 14176
rect 27756 14112 27772 14176
rect 27836 14112 27852 14176
rect 27916 14112 27924 14176
rect 27604 13954 27924 14112
rect 27604 13718 27646 13954
rect 27882 13718 27924 13954
rect 27604 13088 27924 13718
rect 27604 13024 27612 13088
rect 27676 13024 27692 13088
rect 27756 13024 27772 13088
rect 27836 13024 27852 13088
rect 27916 13024 27924 13088
rect 27604 12000 27924 13024
rect 27604 11936 27612 12000
rect 27676 11936 27692 12000
rect 27756 11936 27772 12000
rect 27836 11936 27852 12000
rect 27916 11936 27924 12000
rect 27604 10912 27924 11936
rect 27604 10848 27612 10912
rect 27676 10848 27692 10912
rect 27756 10848 27772 10912
rect 27836 10848 27852 10912
rect 27916 10848 27924 10912
rect 27604 9824 27924 10848
rect 27604 9760 27612 9824
rect 27676 9760 27692 9824
rect 27756 9760 27772 9824
rect 27836 9760 27852 9824
rect 27916 9760 27924 9824
rect 27604 8954 27924 9760
rect 27604 8736 27646 8954
rect 27882 8736 27924 8954
rect 27604 8672 27612 8736
rect 27676 8672 27692 8718
rect 27756 8672 27772 8718
rect 27836 8672 27852 8718
rect 27916 8672 27924 8736
rect 27604 7648 27924 8672
rect 27604 7584 27612 7648
rect 27676 7584 27692 7648
rect 27756 7584 27772 7648
rect 27836 7584 27852 7648
rect 27916 7584 27924 7648
rect 27604 6560 27924 7584
rect 27604 6496 27612 6560
rect 27676 6496 27692 6560
rect 27756 6496 27772 6560
rect 27836 6496 27852 6560
rect 27916 6496 27924 6560
rect 27604 5472 27924 6496
rect 27604 5408 27612 5472
rect 27676 5408 27692 5472
rect 27756 5408 27772 5472
rect 27836 5408 27852 5472
rect 27916 5408 27924 5472
rect 27604 4384 27924 5408
rect 27604 4320 27612 4384
rect 27676 4320 27692 4384
rect 27756 4320 27772 4384
rect 27836 4320 27852 4384
rect 27916 4320 27924 4384
rect 27604 3954 27924 4320
rect 27604 3718 27646 3954
rect 27882 3718 27924 3954
rect 27604 3296 27924 3718
rect 27604 3232 27612 3296
rect 27676 3232 27692 3296
rect 27756 3232 27772 3296
rect 27836 3232 27852 3296
rect 27916 3232 27924 3296
rect 27604 2208 27924 3232
rect 27604 2144 27612 2208
rect 27676 2144 27692 2208
rect 27756 2144 27772 2208
rect 27836 2144 27852 2208
rect 27916 2144 27924 2208
rect 27604 2128 27924 2144
rect 31944 37568 32264 37584
rect 31944 37504 31952 37568
rect 32016 37504 32032 37568
rect 32096 37504 32112 37568
rect 32176 37504 32192 37568
rect 32256 37504 32264 37568
rect 31944 36480 32264 37504
rect 31944 36416 31952 36480
rect 32016 36416 32032 36480
rect 32096 36416 32112 36480
rect 32176 36416 32192 36480
rect 32256 36416 32264 36480
rect 31944 35392 32264 36416
rect 31944 35328 31952 35392
rect 32016 35328 32032 35392
rect 32096 35328 32112 35392
rect 32176 35328 32192 35392
rect 32256 35328 32264 35392
rect 31944 34304 32264 35328
rect 31944 34240 31952 34304
rect 32016 34240 32032 34304
rect 32096 34240 32112 34304
rect 32176 34240 32192 34304
rect 32256 34240 32264 34304
rect 31944 33294 32264 34240
rect 31944 33216 31986 33294
rect 32222 33216 32264 33294
rect 31944 33152 31952 33216
rect 32256 33152 32264 33216
rect 31944 33058 31986 33152
rect 32222 33058 32264 33152
rect 31944 32128 32264 33058
rect 31944 32064 31952 32128
rect 32016 32064 32032 32128
rect 32096 32064 32112 32128
rect 32176 32064 32192 32128
rect 32256 32064 32264 32128
rect 31944 31040 32264 32064
rect 31944 30976 31952 31040
rect 32016 30976 32032 31040
rect 32096 30976 32112 31040
rect 32176 30976 32192 31040
rect 32256 30976 32264 31040
rect 31944 29952 32264 30976
rect 31944 29888 31952 29952
rect 32016 29888 32032 29952
rect 32096 29888 32112 29952
rect 32176 29888 32192 29952
rect 32256 29888 32264 29952
rect 31944 28864 32264 29888
rect 31944 28800 31952 28864
rect 32016 28800 32032 28864
rect 32096 28800 32112 28864
rect 32176 28800 32192 28864
rect 32256 28800 32264 28864
rect 31944 28294 32264 28800
rect 31944 28058 31986 28294
rect 32222 28058 32264 28294
rect 31944 27776 32264 28058
rect 31944 27712 31952 27776
rect 32016 27712 32032 27776
rect 32096 27712 32112 27776
rect 32176 27712 32192 27776
rect 32256 27712 32264 27776
rect 31944 26688 32264 27712
rect 31944 26624 31952 26688
rect 32016 26624 32032 26688
rect 32096 26624 32112 26688
rect 32176 26624 32192 26688
rect 32256 26624 32264 26688
rect 31944 25600 32264 26624
rect 31944 25536 31952 25600
rect 32016 25536 32032 25600
rect 32096 25536 32112 25600
rect 32176 25536 32192 25600
rect 32256 25536 32264 25600
rect 31944 24512 32264 25536
rect 31944 24448 31952 24512
rect 32016 24448 32032 24512
rect 32096 24448 32112 24512
rect 32176 24448 32192 24512
rect 32256 24448 32264 24512
rect 31944 23424 32264 24448
rect 31944 23360 31952 23424
rect 32016 23360 32032 23424
rect 32096 23360 32112 23424
rect 32176 23360 32192 23424
rect 32256 23360 32264 23424
rect 31944 23294 32264 23360
rect 31944 23058 31986 23294
rect 32222 23058 32264 23294
rect 31944 22336 32264 23058
rect 31944 22272 31952 22336
rect 32016 22272 32032 22336
rect 32096 22272 32112 22336
rect 32176 22272 32192 22336
rect 32256 22272 32264 22336
rect 31944 21248 32264 22272
rect 31944 21184 31952 21248
rect 32016 21184 32032 21248
rect 32096 21184 32112 21248
rect 32176 21184 32192 21248
rect 32256 21184 32264 21248
rect 31944 20160 32264 21184
rect 31944 20096 31952 20160
rect 32016 20096 32032 20160
rect 32096 20096 32112 20160
rect 32176 20096 32192 20160
rect 32256 20096 32264 20160
rect 31944 19072 32264 20096
rect 31944 19008 31952 19072
rect 32016 19008 32032 19072
rect 32096 19008 32112 19072
rect 32176 19008 32192 19072
rect 32256 19008 32264 19072
rect 31944 18294 32264 19008
rect 31944 18058 31986 18294
rect 32222 18058 32264 18294
rect 31944 17984 32264 18058
rect 31944 17920 31952 17984
rect 32016 17920 32032 17984
rect 32096 17920 32112 17984
rect 32176 17920 32192 17984
rect 32256 17920 32264 17984
rect 31944 16896 32264 17920
rect 31944 16832 31952 16896
rect 32016 16832 32032 16896
rect 32096 16832 32112 16896
rect 32176 16832 32192 16896
rect 32256 16832 32264 16896
rect 31944 15808 32264 16832
rect 31944 15744 31952 15808
rect 32016 15744 32032 15808
rect 32096 15744 32112 15808
rect 32176 15744 32192 15808
rect 32256 15744 32264 15808
rect 31944 14720 32264 15744
rect 31944 14656 31952 14720
rect 32016 14656 32032 14720
rect 32096 14656 32112 14720
rect 32176 14656 32192 14720
rect 32256 14656 32264 14720
rect 31944 13632 32264 14656
rect 31944 13568 31952 13632
rect 32016 13568 32032 13632
rect 32096 13568 32112 13632
rect 32176 13568 32192 13632
rect 32256 13568 32264 13632
rect 31944 13294 32264 13568
rect 31944 13058 31986 13294
rect 32222 13058 32264 13294
rect 31944 12544 32264 13058
rect 31944 12480 31952 12544
rect 32016 12480 32032 12544
rect 32096 12480 32112 12544
rect 32176 12480 32192 12544
rect 32256 12480 32264 12544
rect 31944 11456 32264 12480
rect 31944 11392 31952 11456
rect 32016 11392 32032 11456
rect 32096 11392 32112 11456
rect 32176 11392 32192 11456
rect 32256 11392 32264 11456
rect 31944 10368 32264 11392
rect 31944 10304 31952 10368
rect 32016 10304 32032 10368
rect 32096 10304 32112 10368
rect 32176 10304 32192 10368
rect 32256 10304 32264 10368
rect 31944 9280 32264 10304
rect 31944 9216 31952 9280
rect 32016 9216 32032 9280
rect 32096 9216 32112 9280
rect 32176 9216 32192 9280
rect 32256 9216 32264 9280
rect 31944 8294 32264 9216
rect 31944 8192 31986 8294
rect 32222 8192 32264 8294
rect 31944 8128 31952 8192
rect 32256 8128 32264 8192
rect 31944 8058 31986 8128
rect 32222 8058 32264 8128
rect 31944 7104 32264 8058
rect 31944 7040 31952 7104
rect 32016 7040 32032 7104
rect 32096 7040 32112 7104
rect 32176 7040 32192 7104
rect 32256 7040 32264 7104
rect 31944 6016 32264 7040
rect 31944 5952 31952 6016
rect 32016 5952 32032 6016
rect 32096 5952 32112 6016
rect 32176 5952 32192 6016
rect 32256 5952 32264 6016
rect 31944 4928 32264 5952
rect 31944 4864 31952 4928
rect 32016 4864 32032 4928
rect 32096 4864 32112 4928
rect 32176 4864 32192 4928
rect 32256 4864 32264 4928
rect 31944 3840 32264 4864
rect 31944 3776 31952 3840
rect 32016 3776 32032 3840
rect 32096 3776 32112 3840
rect 32176 3776 32192 3840
rect 32256 3776 32264 3840
rect 31944 3294 32264 3776
rect 31944 3058 31986 3294
rect 32222 3058 32264 3294
rect 31944 2752 32264 3058
rect 31944 2688 31952 2752
rect 32016 2688 32032 2752
rect 32096 2688 32112 2752
rect 32176 2688 32192 2752
rect 32256 2688 32264 2752
rect 31944 2128 32264 2688
rect 32604 37024 32924 37584
rect 32604 36960 32612 37024
rect 32676 36960 32692 37024
rect 32756 36960 32772 37024
rect 32836 36960 32852 37024
rect 32916 36960 32924 37024
rect 32604 35936 32924 36960
rect 32604 35872 32612 35936
rect 32676 35872 32692 35936
rect 32756 35872 32772 35936
rect 32836 35872 32852 35936
rect 32916 35872 32924 35936
rect 32604 34848 32924 35872
rect 32604 34784 32612 34848
rect 32676 34784 32692 34848
rect 32756 34784 32772 34848
rect 32836 34784 32852 34848
rect 32916 34784 32924 34848
rect 32604 33954 32924 34784
rect 32604 33760 32646 33954
rect 32882 33760 32924 33954
rect 32604 33696 32612 33760
rect 32676 33696 32692 33718
rect 32756 33696 32772 33718
rect 32836 33696 32852 33718
rect 32916 33696 32924 33760
rect 32604 32672 32924 33696
rect 32604 32608 32612 32672
rect 32676 32608 32692 32672
rect 32756 32608 32772 32672
rect 32836 32608 32852 32672
rect 32916 32608 32924 32672
rect 32604 31584 32924 32608
rect 32604 31520 32612 31584
rect 32676 31520 32692 31584
rect 32756 31520 32772 31584
rect 32836 31520 32852 31584
rect 32916 31520 32924 31584
rect 32604 30496 32924 31520
rect 32604 30432 32612 30496
rect 32676 30432 32692 30496
rect 32756 30432 32772 30496
rect 32836 30432 32852 30496
rect 32916 30432 32924 30496
rect 32604 29408 32924 30432
rect 32604 29344 32612 29408
rect 32676 29344 32692 29408
rect 32756 29344 32772 29408
rect 32836 29344 32852 29408
rect 32916 29344 32924 29408
rect 32604 28954 32924 29344
rect 32604 28718 32646 28954
rect 32882 28718 32924 28954
rect 32604 28320 32924 28718
rect 32604 28256 32612 28320
rect 32676 28256 32692 28320
rect 32756 28256 32772 28320
rect 32836 28256 32852 28320
rect 32916 28256 32924 28320
rect 32604 27232 32924 28256
rect 32604 27168 32612 27232
rect 32676 27168 32692 27232
rect 32756 27168 32772 27232
rect 32836 27168 32852 27232
rect 32916 27168 32924 27232
rect 32604 26144 32924 27168
rect 32604 26080 32612 26144
rect 32676 26080 32692 26144
rect 32756 26080 32772 26144
rect 32836 26080 32852 26144
rect 32916 26080 32924 26144
rect 32604 25056 32924 26080
rect 32604 24992 32612 25056
rect 32676 24992 32692 25056
rect 32756 24992 32772 25056
rect 32836 24992 32852 25056
rect 32916 24992 32924 25056
rect 32604 23968 32924 24992
rect 32604 23904 32612 23968
rect 32676 23954 32692 23968
rect 32756 23954 32772 23968
rect 32836 23954 32852 23968
rect 32916 23904 32924 23968
rect 32604 23718 32646 23904
rect 32882 23718 32924 23904
rect 32604 22880 32924 23718
rect 32604 22816 32612 22880
rect 32676 22816 32692 22880
rect 32756 22816 32772 22880
rect 32836 22816 32852 22880
rect 32916 22816 32924 22880
rect 32604 21792 32924 22816
rect 32604 21728 32612 21792
rect 32676 21728 32692 21792
rect 32756 21728 32772 21792
rect 32836 21728 32852 21792
rect 32916 21728 32924 21792
rect 32604 20704 32924 21728
rect 32604 20640 32612 20704
rect 32676 20640 32692 20704
rect 32756 20640 32772 20704
rect 32836 20640 32852 20704
rect 32916 20640 32924 20704
rect 32604 19616 32924 20640
rect 32604 19552 32612 19616
rect 32676 19552 32692 19616
rect 32756 19552 32772 19616
rect 32836 19552 32852 19616
rect 32916 19552 32924 19616
rect 32604 18954 32924 19552
rect 32604 18718 32646 18954
rect 32882 18718 32924 18954
rect 32604 18528 32924 18718
rect 32604 18464 32612 18528
rect 32676 18464 32692 18528
rect 32756 18464 32772 18528
rect 32836 18464 32852 18528
rect 32916 18464 32924 18528
rect 32604 17440 32924 18464
rect 32604 17376 32612 17440
rect 32676 17376 32692 17440
rect 32756 17376 32772 17440
rect 32836 17376 32852 17440
rect 32916 17376 32924 17440
rect 32604 16352 32924 17376
rect 32604 16288 32612 16352
rect 32676 16288 32692 16352
rect 32756 16288 32772 16352
rect 32836 16288 32852 16352
rect 32916 16288 32924 16352
rect 32604 15264 32924 16288
rect 32604 15200 32612 15264
rect 32676 15200 32692 15264
rect 32756 15200 32772 15264
rect 32836 15200 32852 15264
rect 32916 15200 32924 15264
rect 32604 14176 32924 15200
rect 32604 14112 32612 14176
rect 32676 14112 32692 14176
rect 32756 14112 32772 14176
rect 32836 14112 32852 14176
rect 32916 14112 32924 14176
rect 32604 13954 32924 14112
rect 32604 13718 32646 13954
rect 32882 13718 32924 13954
rect 32604 13088 32924 13718
rect 32604 13024 32612 13088
rect 32676 13024 32692 13088
rect 32756 13024 32772 13088
rect 32836 13024 32852 13088
rect 32916 13024 32924 13088
rect 32604 12000 32924 13024
rect 32604 11936 32612 12000
rect 32676 11936 32692 12000
rect 32756 11936 32772 12000
rect 32836 11936 32852 12000
rect 32916 11936 32924 12000
rect 32604 10912 32924 11936
rect 32604 10848 32612 10912
rect 32676 10848 32692 10912
rect 32756 10848 32772 10912
rect 32836 10848 32852 10912
rect 32916 10848 32924 10912
rect 32604 9824 32924 10848
rect 32604 9760 32612 9824
rect 32676 9760 32692 9824
rect 32756 9760 32772 9824
rect 32836 9760 32852 9824
rect 32916 9760 32924 9824
rect 32604 8954 32924 9760
rect 32604 8736 32646 8954
rect 32882 8736 32924 8954
rect 32604 8672 32612 8736
rect 32676 8672 32692 8718
rect 32756 8672 32772 8718
rect 32836 8672 32852 8718
rect 32916 8672 32924 8736
rect 32604 7648 32924 8672
rect 32604 7584 32612 7648
rect 32676 7584 32692 7648
rect 32756 7584 32772 7648
rect 32836 7584 32852 7648
rect 32916 7584 32924 7648
rect 32604 6560 32924 7584
rect 32604 6496 32612 6560
rect 32676 6496 32692 6560
rect 32756 6496 32772 6560
rect 32836 6496 32852 6560
rect 32916 6496 32924 6560
rect 32604 5472 32924 6496
rect 32604 5408 32612 5472
rect 32676 5408 32692 5472
rect 32756 5408 32772 5472
rect 32836 5408 32852 5472
rect 32916 5408 32924 5472
rect 32604 4384 32924 5408
rect 32604 4320 32612 4384
rect 32676 4320 32692 4384
rect 32756 4320 32772 4384
rect 32836 4320 32852 4384
rect 32916 4320 32924 4384
rect 32604 3954 32924 4320
rect 32604 3718 32646 3954
rect 32882 3718 32924 3954
rect 32604 3296 32924 3718
rect 32604 3232 32612 3296
rect 32676 3232 32692 3296
rect 32756 3232 32772 3296
rect 32836 3232 32852 3296
rect 32916 3232 32924 3296
rect 32604 2208 32924 3232
rect 32604 2144 32612 2208
rect 32676 2144 32692 2208
rect 32756 2144 32772 2208
rect 32836 2144 32852 2208
rect 32916 2144 32924 2208
rect 32604 2128 32924 2144
rect 36944 37568 37264 37584
rect 36944 37504 36952 37568
rect 37016 37504 37032 37568
rect 37096 37504 37112 37568
rect 37176 37504 37192 37568
rect 37256 37504 37264 37568
rect 36944 36480 37264 37504
rect 36944 36416 36952 36480
rect 37016 36416 37032 36480
rect 37096 36416 37112 36480
rect 37176 36416 37192 36480
rect 37256 36416 37264 36480
rect 36944 35392 37264 36416
rect 36944 35328 36952 35392
rect 37016 35328 37032 35392
rect 37096 35328 37112 35392
rect 37176 35328 37192 35392
rect 37256 35328 37264 35392
rect 36944 34304 37264 35328
rect 36944 34240 36952 34304
rect 37016 34240 37032 34304
rect 37096 34240 37112 34304
rect 37176 34240 37192 34304
rect 37256 34240 37264 34304
rect 36944 33294 37264 34240
rect 36944 33216 36986 33294
rect 37222 33216 37264 33294
rect 36944 33152 36952 33216
rect 37256 33152 37264 33216
rect 36944 33058 36986 33152
rect 37222 33058 37264 33152
rect 36944 32128 37264 33058
rect 36944 32064 36952 32128
rect 37016 32064 37032 32128
rect 37096 32064 37112 32128
rect 37176 32064 37192 32128
rect 37256 32064 37264 32128
rect 36944 31040 37264 32064
rect 36944 30976 36952 31040
rect 37016 30976 37032 31040
rect 37096 30976 37112 31040
rect 37176 30976 37192 31040
rect 37256 30976 37264 31040
rect 36944 29952 37264 30976
rect 36944 29888 36952 29952
rect 37016 29888 37032 29952
rect 37096 29888 37112 29952
rect 37176 29888 37192 29952
rect 37256 29888 37264 29952
rect 36944 28864 37264 29888
rect 36944 28800 36952 28864
rect 37016 28800 37032 28864
rect 37096 28800 37112 28864
rect 37176 28800 37192 28864
rect 37256 28800 37264 28864
rect 36944 28294 37264 28800
rect 36944 28058 36986 28294
rect 37222 28058 37264 28294
rect 36944 27776 37264 28058
rect 36944 27712 36952 27776
rect 37016 27712 37032 27776
rect 37096 27712 37112 27776
rect 37176 27712 37192 27776
rect 37256 27712 37264 27776
rect 36944 26688 37264 27712
rect 36944 26624 36952 26688
rect 37016 26624 37032 26688
rect 37096 26624 37112 26688
rect 37176 26624 37192 26688
rect 37256 26624 37264 26688
rect 36944 25600 37264 26624
rect 36944 25536 36952 25600
rect 37016 25536 37032 25600
rect 37096 25536 37112 25600
rect 37176 25536 37192 25600
rect 37256 25536 37264 25600
rect 36944 24512 37264 25536
rect 36944 24448 36952 24512
rect 37016 24448 37032 24512
rect 37096 24448 37112 24512
rect 37176 24448 37192 24512
rect 37256 24448 37264 24512
rect 36944 23424 37264 24448
rect 36944 23360 36952 23424
rect 37016 23360 37032 23424
rect 37096 23360 37112 23424
rect 37176 23360 37192 23424
rect 37256 23360 37264 23424
rect 36944 23294 37264 23360
rect 36944 23058 36986 23294
rect 37222 23058 37264 23294
rect 36944 22336 37264 23058
rect 36944 22272 36952 22336
rect 37016 22272 37032 22336
rect 37096 22272 37112 22336
rect 37176 22272 37192 22336
rect 37256 22272 37264 22336
rect 36944 21248 37264 22272
rect 36944 21184 36952 21248
rect 37016 21184 37032 21248
rect 37096 21184 37112 21248
rect 37176 21184 37192 21248
rect 37256 21184 37264 21248
rect 36944 20160 37264 21184
rect 36944 20096 36952 20160
rect 37016 20096 37032 20160
rect 37096 20096 37112 20160
rect 37176 20096 37192 20160
rect 37256 20096 37264 20160
rect 36944 19072 37264 20096
rect 36944 19008 36952 19072
rect 37016 19008 37032 19072
rect 37096 19008 37112 19072
rect 37176 19008 37192 19072
rect 37256 19008 37264 19072
rect 36944 18294 37264 19008
rect 36944 18058 36986 18294
rect 37222 18058 37264 18294
rect 36944 17984 37264 18058
rect 36944 17920 36952 17984
rect 37016 17920 37032 17984
rect 37096 17920 37112 17984
rect 37176 17920 37192 17984
rect 37256 17920 37264 17984
rect 36944 16896 37264 17920
rect 36944 16832 36952 16896
rect 37016 16832 37032 16896
rect 37096 16832 37112 16896
rect 37176 16832 37192 16896
rect 37256 16832 37264 16896
rect 36944 15808 37264 16832
rect 36944 15744 36952 15808
rect 37016 15744 37032 15808
rect 37096 15744 37112 15808
rect 37176 15744 37192 15808
rect 37256 15744 37264 15808
rect 36944 14720 37264 15744
rect 36944 14656 36952 14720
rect 37016 14656 37032 14720
rect 37096 14656 37112 14720
rect 37176 14656 37192 14720
rect 37256 14656 37264 14720
rect 36944 13632 37264 14656
rect 36944 13568 36952 13632
rect 37016 13568 37032 13632
rect 37096 13568 37112 13632
rect 37176 13568 37192 13632
rect 37256 13568 37264 13632
rect 36944 13294 37264 13568
rect 36944 13058 36986 13294
rect 37222 13058 37264 13294
rect 36944 12544 37264 13058
rect 36944 12480 36952 12544
rect 37016 12480 37032 12544
rect 37096 12480 37112 12544
rect 37176 12480 37192 12544
rect 37256 12480 37264 12544
rect 36944 11456 37264 12480
rect 36944 11392 36952 11456
rect 37016 11392 37032 11456
rect 37096 11392 37112 11456
rect 37176 11392 37192 11456
rect 37256 11392 37264 11456
rect 36944 10368 37264 11392
rect 36944 10304 36952 10368
rect 37016 10304 37032 10368
rect 37096 10304 37112 10368
rect 37176 10304 37192 10368
rect 37256 10304 37264 10368
rect 36944 9280 37264 10304
rect 36944 9216 36952 9280
rect 37016 9216 37032 9280
rect 37096 9216 37112 9280
rect 37176 9216 37192 9280
rect 37256 9216 37264 9280
rect 36944 8294 37264 9216
rect 36944 8192 36986 8294
rect 37222 8192 37264 8294
rect 36944 8128 36952 8192
rect 37256 8128 37264 8192
rect 36944 8058 36986 8128
rect 37222 8058 37264 8128
rect 36944 7104 37264 8058
rect 36944 7040 36952 7104
rect 37016 7040 37032 7104
rect 37096 7040 37112 7104
rect 37176 7040 37192 7104
rect 37256 7040 37264 7104
rect 36944 6016 37264 7040
rect 36944 5952 36952 6016
rect 37016 5952 37032 6016
rect 37096 5952 37112 6016
rect 37176 5952 37192 6016
rect 37256 5952 37264 6016
rect 36944 4928 37264 5952
rect 36944 4864 36952 4928
rect 37016 4864 37032 4928
rect 37096 4864 37112 4928
rect 37176 4864 37192 4928
rect 37256 4864 37264 4928
rect 36944 3840 37264 4864
rect 36944 3776 36952 3840
rect 37016 3776 37032 3840
rect 37096 3776 37112 3840
rect 37176 3776 37192 3840
rect 37256 3776 37264 3840
rect 36944 3294 37264 3776
rect 36944 3058 36986 3294
rect 37222 3058 37264 3294
rect 36944 2752 37264 3058
rect 36944 2688 36952 2752
rect 37016 2688 37032 2752
rect 37096 2688 37112 2752
rect 37176 2688 37192 2752
rect 37256 2688 37264 2752
rect 36944 2128 37264 2688
rect 37604 37024 37924 37584
rect 37604 36960 37612 37024
rect 37676 36960 37692 37024
rect 37756 36960 37772 37024
rect 37836 36960 37852 37024
rect 37916 36960 37924 37024
rect 37604 35936 37924 36960
rect 37604 35872 37612 35936
rect 37676 35872 37692 35936
rect 37756 35872 37772 35936
rect 37836 35872 37852 35936
rect 37916 35872 37924 35936
rect 37604 34848 37924 35872
rect 37604 34784 37612 34848
rect 37676 34784 37692 34848
rect 37756 34784 37772 34848
rect 37836 34784 37852 34848
rect 37916 34784 37924 34848
rect 37604 33954 37924 34784
rect 37604 33760 37646 33954
rect 37882 33760 37924 33954
rect 37604 33696 37612 33760
rect 37676 33696 37692 33718
rect 37756 33696 37772 33718
rect 37836 33696 37852 33718
rect 37916 33696 37924 33760
rect 37604 32672 37924 33696
rect 37604 32608 37612 32672
rect 37676 32608 37692 32672
rect 37756 32608 37772 32672
rect 37836 32608 37852 32672
rect 37916 32608 37924 32672
rect 37604 31584 37924 32608
rect 37604 31520 37612 31584
rect 37676 31520 37692 31584
rect 37756 31520 37772 31584
rect 37836 31520 37852 31584
rect 37916 31520 37924 31584
rect 37604 30496 37924 31520
rect 37604 30432 37612 30496
rect 37676 30432 37692 30496
rect 37756 30432 37772 30496
rect 37836 30432 37852 30496
rect 37916 30432 37924 30496
rect 37604 29408 37924 30432
rect 37604 29344 37612 29408
rect 37676 29344 37692 29408
rect 37756 29344 37772 29408
rect 37836 29344 37852 29408
rect 37916 29344 37924 29408
rect 37604 28954 37924 29344
rect 37604 28718 37646 28954
rect 37882 28718 37924 28954
rect 37604 28320 37924 28718
rect 37604 28256 37612 28320
rect 37676 28256 37692 28320
rect 37756 28256 37772 28320
rect 37836 28256 37852 28320
rect 37916 28256 37924 28320
rect 37604 27232 37924 28256
rect 37604 27168 37612 27232
rect 37676 27168 37692 27232
rect 37756 27168 37772 27232
rect 37836 27168 37852 27232
rect 37916 27168 37924 27232
rect 37604 26144 37924 27168
rect 37604 26080 37612 26144
rect 37676 26080 37692 26144
rect 37756 26080 37772 26144
rect 37836 26080 37852 26144
rect 37916 26080 37924 26144
rect 37604 25056 37924 26080
rect 37604 24992 37612 25056
rect 37676 24992 37692 25056
rect 37756 24992 37772 25056
rect 37836 24992 37852 25056
rect 37916 24992 37924 25056
rect 37604 23968 37924 24992
rect 37604 23904 37612 23968
rect 37676 23954 37692 23968
rect 37756 23954 37772 23968
rect 37836 23954 37852 23968
rect 37916 23904 37924 23968
rect 37604 23718 37646 23904
rect 37882 23718 37924 23904
rect 37604 22880 37924 23718
rect 37604 22816 37612 22880
rect 37676 22816 37692 22880
rect 37756 22816 37772 22880
rect 37836 22816 37852 22880
rect 37916 22816 37924 22880
rect 37604 21792 37924 22816
rect 37604 21728 37612 21792
rect 37676 21728 37692 21792
rect 37756 21728 37772 21792
rect 37836 21728 37852 21792
rect 37916 21728 37924 21792
rect 37604 20704 37924 21728
rect 37604 20640 37612 20704
rect 37676 20640 37692 20704
rect 37756 20640 37772 20704
rect 37836 20640 37852 20704
rect 37916 20640 37924 20704
rect 37604 19616 37924 20640
rect 37604 19552 37612 19616
rect 37676 19552 37692 19616
rect 37756 19552 37772 19616
rect 37836 19552 37852 19616
rect 37916 19552 37924 19616
rect 37604 18954 37924 19552
rect 37604 18718 37646 18954
rect 37882 18718 37924 18954
rect 37604 18528 37924 18718
rect 37604 18464 37612 18528
rect 37676 18464 37692 18528
rect 37756 18464 37772 18528
rect 37836 18464 37852 18528
rect 37916 18464 37924 18528
rect 37604 17440 37924 18464
rect 37604 17376 37612 17440
rect 37676 17376 37692 17440
rect 37756 17376 37772 17440
rect 37836 17376 37852 17440
rect 37916 17376 37924 17440
rect 37604 16352 37924 17376
rect 37604 16288 37612 16352
rect 37676 16288 37692 16352
rect 37756 16288 37772 16352
rect 37836 16288 37852 16352
rect 37916 16288 37924 16352
rect 37604 15264 37924 16288
rect 37604 15200 37612 15264
rect 37676 15200 37692 15264
rect 37756 15200 37772 15264
rect 37836 15200 37852 15264
rect 37916 15200 37924 15264
rect 37604 14176 37924 15200
rect 37604 14112 37612 14176
rect 37676 14112 37692 14176
rect 37756 14112 37772 14176
rect 37836 14112 37852 14176
rect 37916 14112 37924 14176
rect 37604 13954 37924 14112
rect 37604 13718 37646 13954
rect 37882 13718 37924 13954
rect 37604 13088 37924 13718
rect 37604 13024 37612 13088
rect 37676 13024 37692 13088
rect 37756 13024 37772 13088
rect 37836 13024 37852 13088
rect 37916 13024 37924 13088
rect 37604 12000 37924 13024
rect 37604 11936 37612 12000
rect 37676 11936 37692 12000
rect 37756 11936 37772 12000
rect 37836 11936 37852 12000
rect 37916 11936 37924 12000
rect 37604 10912 37924 11936
rect 37604 10848 37612 10912
rect 37676 10848 37692 10912
rect 37756 10848 37772 10912
rect 37836 10848 37852 10912
rect 37916 10848 37924 10912
rect 37604 9824 37924 10848
rect 37604 9760 37612 9824
rect 37676 9760 37692 9824
rect 37756 9760 37772 9824
rect 37836 9760 37852 9824
rect 37916 9760 37924 9824
rect 37604 8954 37924 9760
rect 37604 8736 37646 8954
rect 37882 8736 37924 8954
rect 37604 8672 37612 8736
rect 37676 8672 37692 8718
rect 37756 8672 37772 8718
rect 37836 8672 37852 8718
rect 37916 8672 37924 8736
rect 37604 7648 37924 8672
rect 37604 7584 37612 7648
rect 37676 7584 37692 7648
rect 37756 7584 37772 7648
rect 37836 7584 37852 7648
rect 37916 7584 37924 7648
rect 37604 6560 37924 7584
rect 37604 6496 37612 6560
rect 37676 6496 37692 6560
rect 37756 6496 37772 6560
rect 37836 6496 37852 6560
rect 37916 6496 37924 6560
rect 37604 5472 37924 6496
rect 37604 5408 37612 5472
rect 37676 5408 37692 5472
rect 37756 5408 37772 5472
rect 37836 5408 37852 5472
rect 37916 5408 37924 5472
rect 37604 4384 37924 5408
rect 37604 4320 37612 4384
rect 37676 4320 37692 4384
rect 37756 4320 37772 4384
rect 37836 4320 37852 4384
rect 37916 4320 37924 4384
rect 37604 3954 37924 4320
rect 37604 3718 37646 3954
rect 37882 3718 37924 3954
rect 37604 3296 37924 3718
rect 37604 3232 37612 3296
rect 37676 3232 37692 3296
rect 37756 3232 37772 3296
rect 37836 3232 37852 3296
rect 37916 3232 37924 3296
rect 37604 2208 37924 3232
rect 37604 2144 37612 2208
rect 37676 2144 37692 2208
rect 37756 2144 37772 2208
rect 37836 2144 37852 2208
rect 37916 2144 37924 2208
rect 37604 2128 37924 2144
<< via4 >>
rect 1986 33216 2222 33294
rect 1986 33152 2016 33216
rect 2016 33152 2032 33216
rect 2032 33152 2096 33216
rect 2096 33152 2112 33216
rect 2112 33152 2176 33216
rect 2176 33152 2192 33216
rect 2192 33152 2222 33216
rect 1986 33058 2222 33152
rect 1986 28058 2222 28294
rect 1986 23058 2222 23294
rect 1986 18058 2222 18294
rect 1986 13058 2222 13294
rect 1986 8192 2222 8294
rect 1986 8128 2016 8192
rect 2016 8128 2032 8192
rect 2032 8128 2096 8192
rect 2096 8128 2112 8192
rect 2112 8128 2176 8192
rect 2176 8128 2192 8192
rect 2192 8128 2222 8192
rect 1986 8058 2222 8128
rect 1986 3058 2222 3294
rect 2646 33760 2882 33954
rect 2646 33718 2676 33760
rect 2676 33718 2692 33760
rect 2692 33718 2756 33760
rect 2756 33718 2772 33760
rect 2772 33718 2836 33760
rect 2836 33718 2852 33760
rect 2852 33718 2882 33760
rect 2646 28718 2882 28954
rect 2646 23904 2676 23954
rect 2676 23904 2692 23954
rect 2692 23904 2756 23954
rect 2756 23904 2772 23954
rect 2772 23904 2836 23954
rect 2836 23904 2852 23954
rect 2852 23904 2882 23954
rect 2646 23718 2882 23904
rect 2646 18718 2882 18954
rect 2646 13718 2882 13954
rect 2646 8736 2882 8954
rect 2646 8718 2676 8736
rect 2676 8718 2692 8736
rect 2692 8718 2756 8736
rect 2756 8718 2772 8736
rect 2772 8718 2836 8736
rect 2836 8718 2852 8736
rect 2852 8718 2882 8736
rect 2646 3718 2882 3954
rect 6986 33216 7222 33294
rect 6986 33152 7016 33216
rect 7016 33152 7032 33216
rect 7032 33152 7096 33216
rect 7096 33152 7112 33216
rect 7112 33152 7176 33216
rect 7176 33152 7192 33216
rect 7192 33152 7222 33216
rect 6986 33058 7222 33152
rect 6986 28058 7222 28294
rect 6986 23058 7222 23294
rect 6986 18058 7222 18294
rect 6986 13058 7222 13294
rect 6986 8192 7222 8294
rect 6986 8128 7016 8192
rect 7016 8128 7032 8192
rect 7032 8128 7096 8192
rect 7096 8128 7112 8192
rect 7112 8128 7176 8192
rect 7176 8128 7192 8192
rect 7192 8128 7222 8192
rect 6986 8058 7222 8128
rect 6986 3058 7222 3294
rect 7646 33760 7882 33954
rect 7646 33718 7676 33760
rect 7676 33718 7692 33760
rect 7692 33718 7756 33760
rect 7756 33718 7772 33760
rect 7772 33718 7836 33760
rect 7836 33718 7852 33760
rect 7852 33718 7882 33760
rect 7646 28718 7882 28954
rect 7646 23904 7676 23954
rect 7676 23904 7692 23954
rect 7692 23904 7756 23954
rect 7756 23904 7772 23954
rect 7772 23904 7836 23954
rect 7836 23904 7852 23954
rect 7852 23904 7882 23954
rect 7646 23718 7882 23904
rect 7646 18718 7882 18954
rect 7646 13718 7882 13954
rect 7646 8736 7882 8954
rect 7646 8718 7676 8736
rect 7676 8718 7692 8736
rect 7692 8718 7756 8736
rect 7756 8718 7772 8736
rect 7772 8718 7836 8736
rect 7836 8718 7852 8736
rect 7852 8718 7882 8736
rect 7646 3718 7882 3954
rect 11986 33216 12222 33294
rect 11986 33152 12016 33216
rect 12016 33152 12032 33216
rect 12032 33152 12096 33216
rect 12096 33152 12112 33216
rect 12112 33152 12176 33216
rect 12176 33152 12192 33216
rect 12192 33152 12222 33216
rect 11986 33058 12222 33152
rect 11986 28058 12222 28294
rect 11986 23058 12222 23294
rect 11986 18058 12222 18294
rect 11986 13058 12222 13294
rect 11986 8192 12222 8294
rect 11986 8128 12016 8192
rect 12016 8128 12032 8192
rect 12032 8128 12096 8192
rect 12096 8128 12112 8192
rect 12112 8128 12176 8192
rect 12176 8128 12192 8192
rect 12192 8128 12222 8192
rect 11986 8058 12222 8128
rect 11986 3058 12222 3294
rect 12646 33760 12882 33954
rect 12646 33718 12676 33760
rect 12676 33718 12692 33760
rect 12692 33718 12756 33760
rect 12756 33718 12772 33760
rect 12772 33718 12836 33760
rect 12836 33718 12852 33760
rect 12852 33718 12882 33760
rect 12646 28718 12882 28954
rect 12646 23904 12676 23954
rect 12676 23904 12692 23954
rect 12692 23904 12756 23954
rect 12756 23904 12772 23954
rect 12772 23904 12836 23954
rect 12836 23904 12852 23954
rect 12852 23904 12882 23954
rect 12646 23718 12882 23904
rect 12646 18718 12882 18954
rect 12646 13718 12882 13954
rect 12646 8736 12882 8954
rect 12646 8718 12676 8736
rect 12676 8718 12692 8736
rect 12692 8718 12756 8736
rect 12756 8718 12772 8736
rect 12772 8718 12836 8736
rect 12836 8718 12852 8736
rect 12852 8718 12882 8736
rect 12646 3718 12882 3954
rect 16986 33216 17222 33294
rect 16986 33152 17016 33216
rect 17016 33152 17032 33216
rect 17032 33152 17096 33216
rect 17096 33152 17112 33216
rect 17112 33152 17176 33216
rect 17176 33152 17192 33216
rect 17192 33152 17222 33216
rect 16986 33058 17222 33152
rect 16986 28058 17222 28294
rect 16986 23058 17222 23294
rect 16986 18058 17222 18294
rect 16986 13058 17222 13294
rect 16986 8192 17222 8294
rect 16986 8128 17016 8192
rect 17016 8128 17032 8192
rect 17032 8128 17096 8192
rect 17096 8128 17112 8192
rect 17112 8128 17176 8192
rect 17176 8128 17192 8192
rect 17192 8128 17222 8192
rect 16986 8058 17222 8128
rect 16986 3058 17222 3294
rect 17646 33760 17882 33954
rect 17646 33718 17676 33760
rect 17676 33718 17692 33760
rect 17692 33718 17756 33760
rect 17756 33718 17772 33760
rect 17772 33718 17836 33760
rect 17836 33718 17852 33760
rect 17852 33718 17882 33760
rect 17646 28718 17882 28954
rect 17646 23904 17676 23954
rect 17676 23904 17692 23954
rect 17692 23904 17756 23954
rect 17756 23904 17772 23954
rect 17772 23904 17836 23954
rect 17836 23904 17852 23954
rect 17852 23904 17882 23954
rect 17646 23718 17882 23904
rect 17646 18718 17882 18954
rect 17646 13718 17882 13954
rect 17646 8736 17882 8954
rect 17646 8718 17676 8736
rect 17676 8718 17692 8736
rect 17692 8718 17756 8736
rect 17756 8718 17772 8736
rect 17772 8718 17836 8736
rect 17836 8718 17852 8736
rect 17852 8718 17882 8736
rect 17646 3718 17882 3954
rect 21986 33216 22222 33294
rect 21986 33152 22016 33216
rect 22016 33152 22032 33216
rect 22032 33152 22096 33216
rect 22096 33152 22112 33216
rect 22112 33152 22176 33216
rect 22176 33152 22192 33216
rect 22192 33152 22222 33216
rect 21986 33058 22222 33152
rect 21986 28058 22222 28294
rect 21986 23058 22222 23294
rect 21986 18058 22222 18294
rect 21986 13058 22222 13294
rect 21986 8192 22222 8294
rect 21986 8128 22016 8192
rect 22016 8128 22032 8192
rect 22032 8128 22096 8192
rect 22096 8128 22112 8192
rect 22112 8128 22176 8192
rect 22176 8128 22192 8192
rect 22192 8128 22222 8192
rect 21986 8058 22222 8128
rect 21986 3058 22222 3294
rect 22646 33760 22882 33954
rect 22646 33718 22676 33760
rect 22676 33718 22692 33760
rect 22692 33718 22756 33760
rect 22756 33718 22772 33760
rect 22772 33718 22836 33760
rect 22836 33718 22852 33760
rect 22852 33718 22882 33760
rect 22646 28718 22882 28954
rect 22646 23904 22676 23954
rect 22676 23904 22692 23954
rect 22692 23904 22756 23954
rect 22756 23904 22772 23954
rect 22772 23904 22836 23954
rect 22836 23904 22852 23954
rect 22852 23904 22882 23954
rect 22646 23718 22882 23904
rect 22646 18718 22882 18954
rect 22646 13718 22882 13954
rect 22646 8736 22882 8954
rect 22646 8718 22676 8736
rect 22676 8718 22692 8736
rect 22692 8718 22756 8736
rect 22756 8718 22772 8736
rect 22772 8718 22836 8736
rect 22836 8718 22852 8736
rect 22852 8718 22882 8736
rect 22646 3718 22882 3954
rect 26986 33216 27222 33294
rect 26986 33152 27016 33216
rect 27016 33152 27032 33216
rect 27032 33152 27096 33216
rect 27096 33152 27112 33216
rect 27112 33152 27176 33216
rect 27176 33152 27192 33216
rect 27192 33152 27222 33216
rect 26986 33058 27222 33152
rect 26986 28058 27222 28294
rect 26986 23058 27222 23294
rect 26986 18058 27222 18294
rect 26986 13058 27222 13294
rect 26986 8192 27222 8294
rect 26986 8128 27016 8192
rect 27016 8128 27032 8192
rect 27032 8128 27096 8192
rect 27096 8128 27112 8192
rect 27112 8128 27176 8192
rect 27176 8128 27192 8192
rect 27192 8128 27222 8192
rect 26986 8058 27222 8128
rect 26986 3058 27222 3294
rect 27646 33760 27882 33954
rect 27646 33718 27676 33760
rect 27676 33718 27692 33760
rect 27692 33718 27756 33760
rect 27756 33718 27772 33760
rect 27772 33718 27836 33760
rect 27836 33718 27852 33760
rect 27852 33718 27882 33760
rect 27646 28718 27882 28954
rect 27646 23904 27676 23954
rect 27676 23904 27692 23954
rect 27692 23904 27756 23954
rect 27756 23904 27772 23954
rect 27772 23904 27836 23954
rect 27836 23904 27852 23954
rect 27852 23904 27882 23954
rect 27646 23718 27882 23904
rect 27646 18718 27882 18954
rect 27646 13718 27882 13954
rect 27646 8736 27882 8954
rect 27646 8718 27676 8736
rect 27676 8718 27692 8736
rect 27692 8718 27756 8736
rect 27756 8718 27772 8736
rect 27772 8718 27836 8736
rect 27836 8718 27852 8736
rect 27852 8718 27882 8736
rect 27646 3718 27882 3954
rect 31986 33216 32222 33294
rect 31986 33152 32016 33216
rect 32016 33152 32032 33216
rect 32032 33152 32096 33216
rect 32096 33152 32112 33216
rect 32112 33152 32176 33216
rect 32176 33152 32192 33216
rect 32192 33152 32222 33216
rect 31986 33058 32222 33152
rect 31986 28058 32222 28294
rect 31986 23058 32222 23294
rect 31986 18058 32222 18294
rect 31986 13058 32222 13294
rect 31986 8192 32222 8294
rect 31986 8128 32016 8192
rect 32016 8128 32032 8192
rect 32032 8128 32096 8192
rect 32096 8128 32112 8192
rect 32112 8128 32176 8192
rect 32176 8128 32192 8192
rect 32192 8128 32222 8192
rect 31986 8058 32222 8128
rect 31986 3058 32222 3294
rect 32646 33760 32882 33954
rect 32646 33718 32676 33760
rect 32676 33718 32692 33760
rect 32692 33718 32756 33760
rect 32756 33718 32772 33760
rect 32772 33718 32836 33760
rect 32836 33718 32852 33760
rect 32852 33718 32882 33760
rect 32646 28718 32882 28954
rect 32646 23904 32676 23954
rect 32676 23904 32692 23954
rect 32692 23904 32756 23954
rect 32756 23904 32772 23954
rect 32772 23904 32836 23954
rect 32836 23904 32852 23954
rect 32852 23904 32882 23954
rect 32646 23718 32882 23904
rect 32646 18718 32882 18954
rect 32646 13718 32882 13954
rect 32646 8736 32882 8954
rect 32646 8718 32676 8736
rect 32676 8718 32692 8736
rect 32692 8718 32756 8736
rect 32756 8718 32772 8736
rect 32772 8718 32836 8736
rect 32836 8718 32852 8736
rect 32852 8718 32882 8736
rect 32646 3718 32882 3954
rect 36986 33216 37222 33294
rect 36986 33152 37016 33216
rect 37016 33152 37032 33216
rect 37032 33152 37096 33216
rect 37096 33152 37112 33216
rect 37112 33152 37176 33216
rect 37176 33152 37192 33216
rect 37192 33152 37222 33216
rect 36986 33058 37222 33152
rect 36986 28058 37222 28294
rect 36986 23058 37222 23294
rect 36986 18058 37222 18294
rect 36986 13058 37222 13294
rect 36986 8192 37222 8294
rect 36986 8128 37016 8192
rect 37016 8128 37032 8192
rect 37032 8128 37096 8192
rect 37096 8128 37112 8192
rect 37112 8128 37176 8192
rect 37176 8128 37192 8192
rect 37192 8128 37222 8192
rect 36986 8058 37222 8128
rect 36986 3058 37222 3294
rect 37646 33760 37882 33954
rect 37646 33718 37676 33760
rect 37676 33718 37692 33760
rect 37692 33718 37756 33760
rect 37756 33718 37772 33760
rect 37772 33718 37836 33760
rect 37836 33718 37852 33760
rect 37852 33718 37882 33760
rect 37646 28718 37882 28954
rect 37646 23904 37676 23954
rect 37676 23904 37692 23954
rect 37692 23904 37756 23954
rect 37756 23904 37772 23954
rect 37772 23904 37836 23954
rect 37836 23904 37852 23954
rect 37852 23904 37882 23954
rect 37646 23718 37882 23904
rect 37646 18718 37882 18954
rect 37646 13718 37882 13954
rect 37646 8736 37882 8954
rect 37646 8718 37676 8736
rect 37676 8718 37692 8736
rect 37692 8718 37756 8736
rect 37756 8718 37772 8736
rect 37772 8718 37836 8736
rect 37836 8718 37852 8736
rect 37852 8718 37882 8736
rect 37646 3718 37882 3954
<< metal5 >>
rect 1056 33954 38872 33996
rect 1056 33718 2646 33954
rect 2882 33718 7646 33954
rect 7882 33718 12646 33954
rect 12882 33718 17646 33954
rect 17882 33718 22646 33954
rect 22882 33718 27646 33954
rect 27882 33718 32646 33954
rect 32882 33718 37646 33954
rect 37882 33718 38872 33954
rect 1056 33676 38872 33718
rect 1056 33294 38872 33336
rect 1056 33058 1986 33294
rect 2222 33058 6986 33294
rect 7222 33058 11986 33294
rect 12222 33058 16986 33294
rect 17222 33058 21986 33294
rect 22222 33058 26986 33294
rect 27222 33058 31986 33294
rect 32222 33058 36986 33294
rect 37222 33058 38872 33294
rect 1056 33016 38872 33058
rect 1056 28954 38872 28996
rect 1056 28718 2646 28954
rect 2882 28718 7646 28954
rect 7882 28718 12646 28954
rect 12882 28718 17646 28954
rect 17882 28718 22646 28954
rect 22882 28718 27646 28954
rect 27882 28718 32646 28954
rect 32882 28718 37646 28954
rect 37882 28718 38872 28954
rect 1056 28676 38872 28718
rect 1056 28294 38872 28336
rect 1056 28058 1986 28294
rect 2222 28058 6986 28294
rect 7222 28058 11986 28294
rect 12222 28058 16986 28294
rect 17222 28058 21986 28294
rect 22222 28058 26986 28294
rect 27222 28058 31986 28294
rect 32222 28058 36986 28294
rect 37222 28058 38872 28294
rect 1056 28016 38872 28058
rect 1056 23954 38872 23996
rect 1056 23718 2646 23954
rect 2882 23718 7646 23954
rect 7882 23718 12646 23954
rect 12882 23718 17646 23954
rect 17882 23718 22646 23954
rect 22882 23718 27646 23954
rect 27882 23718 32646 23954
rect 32882 23718 37646 23954
rect 37882 23718 38872 23954
rect 1056 23676 38872 23718
rect 1056 23294 38872 23336
rect 1056 23058 1986 23294
rect 2222 23058 6986 23294
rect 7222 23058 11986 23294
rect 12222 23058 16986 23294
rect 17222 23058 21986 23294
rect 22222 23058 26986 23294
rect 27222 23058 31986 23294
rect 32222 23058 36986 23294
rect 37222 23058 38872 23294
rect 1056 23016 38872 23058
rect 1056 18954 38872 18996
rect 1056 18718 2646 18954
rect 2882 18718 7646 18954
rect 7882 18718 12646 18954
rect 12882 18718 17646 18954
rect 17882 18718 22646 18954
rect 22882 18718 27646 18954
rect 27882 18718 32646 18954
rect 32882 18718 37646 18954
rect 37882 18718 38872 18954
rect 1056 18676 38872 18718
rect 1056 18294 38872 18336
rect 1056 18058 1986 18294
rect 2222 18058 6986 18294
rect 7222 18058 11986 18294
rect 12222 18058 16986 18294
rect 17222 18058 21986 18294
rect 22222 18058 26986 18294
rect 27222 18058 31986 18294
rect 32222 18058 36986 18294
rect 37222 18058 38872 18294
rect 1056 18016 38872 18058
rect 1056 13954 38872 13996
rect 1056 13718 2646 13954
rect 2882 13718 7646 13954
rect 7882 13718 12646 13954
rect 12882 13718 17646 13954
rect 17882 13718 22646 13954
rect 22882 13718 27646 13954
rect 27882 13718 32646 13954
rect 32882 13718 37646 13954
rect 37882 13718 38872 13954
rect 1056 13676 38872 13718
rect 1056 13294 38872 13336
rect 1056 13058 1986 13294
rect 2222 13058 6986 13294
rect 7222 13058 11986 13294
rect 12222 13058 16986 13294
rect 17222 13058 21986 13294
rect 22222 13058 26986 13294
rect 27222 13058 31986 13294
rect 32222 13058 36986 13294
rect 37222 13058 38872 13294
rect 1056 13016 38872 13058
rect 1056 8954 38872 8996
rect 1056 8718 2646 8954
rect 2882 8718 7646 8954
rect 7882 8718 12646 8954
rect 12882 8718 17646 8954
rect 17882 8718 22646 8954
rect 22882 8718 27646 8954
rect 27882 8718 32646 8954
rect 32882 8718 37646 8954
rect 37882 8718 38872 8954
rect 1056 8676 38872 8718
rect 1056 8294 38872 8336
rect 1056 8058 1986 8294
rect 2222 8058 6986 8294
rect 7222 8058 11986 8294
rect 12222 8058 16986 8294
rect 17222 8058 21986 8294
rect 22222 8058 26986 8294
rect 27222 8058 31986 8294
rect 32222 8058 36986 8294
rect 37222 8058 38872 8294
rect 1056 8016 38872 8058
rect 1056 3954 38872 3996
rect 1056 3718 2646 3954
rect 2882 3718 7646 3954
rect 7882 3718 12646 3954
rect 12882 3718 17646 3954
rect 17882 3718 22646 3954
rect 22882 3718 27646 3954
rect 27882 3718 32646 3954
rect 32882 3718 37646 3954
rect 37882 3718 38872 3954
rect 1056 3676 38872 3718
rect 1056 3294 38872 3336
rect 1056 3058 1986 3294
rect 2222 3058 6986 3294
rect 7222 3058 11986 3294
rect 12222 3058 16986 3294
rect 17222 3058 21986 3294
rect 22222 3058 26986 3294
rect 27222 3058 31986 3294
rect 32222 3058 36986 3294
rect 37222 3058 38872 3294
rect 1056 3016 38872 3058
use sky130_fd_sc_hd__and4_2  clk_sky130_fd_sc_hd__and4_2_D
timestamp 0
transform 1 0 20424 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_2  clk_sky130_fd_sc_hd__and4b_2_B
timestamp 0
transform 1 0 19504 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_2  clk_sky130_fd_sc_hd__and4b_2_C
timestamp 0
transform 1 0 18308 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_2  clk_sky130_fd_sc_hd__and4b_2_D
timestamp 0
transform 1 0 19504 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_2  clk_sky130_fd_sc_hd__and4bb_2_C_1
timestamp 0
transform 1 0 19504 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_2  clk_sky130_fd_sc_hd__and4bb_2_C
timestamp 0
transform 1 0 19504 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_2  clk_sky130_fd_sc_hd__and4bb_2_D
timestamp 0
transform 1 0 20424 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 21804 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 0
transform -1 0 20516 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 0
transform 1 0 21436 0 1 18496
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 0
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 0
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 0
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 0
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 0
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 0
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 0
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 0
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 0
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 0
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 0
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 0
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 0
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 0
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 0
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 0
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 0
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 0
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 0
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_405
timestamp 0
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 0
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 0
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 0
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 0
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 0
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 0
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 0
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 0
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 0
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 0
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 0
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 0
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 0
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 0
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 0
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 0
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 0
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 0
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 0
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 0
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 0
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 0
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_405
timestamp 0
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 0
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 0
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 0
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 0
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 0
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 0
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 0
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 0
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 0
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 0
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 0
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 0
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 0
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 0
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 0
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 0
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 0
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 0
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 0
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 0
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 0
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 0
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 0
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_401
timestamp 0
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 0
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 0
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 0
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 0
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 0
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 0
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 0
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 0
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 0
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 0
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 0
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 0
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 0
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 0
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 0
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 0
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 0
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 0
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 0
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 0
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 0
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 0
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 0
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 0
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_405
timestamp 0
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 0
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 0
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 0
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 0
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 0
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 0
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 0
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 0
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 0
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 0
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 0
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 0
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 0
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 0
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 0
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 0
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 0
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 0
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 0
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 0
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 0
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 0
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 0
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 0
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 0
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 0
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_401
timestamp 0
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 0
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 0
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 0
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 0
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 0
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 0
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 0
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 0
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 0
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 0
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 0
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 0
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 0
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 0
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 0
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 0
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 0
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 0
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 0
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 0
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 0
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 0
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 0
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 0
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 0
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 0
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_405
timestamp 0
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 0
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 0
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 0
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 0
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 0
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 0
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 0
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 0
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 0
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 0
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 0
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 0
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 0
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 0
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 0
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 0
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 0
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 0
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 0
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 0
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 0
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 0
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 0
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 0
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 0
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 0
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_401
timestamp 0
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 0
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 0
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 0
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 0
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 0
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 0
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 0
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 0
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 0
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 0
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 0
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 0
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 0
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 0
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 0
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 0
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 0
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 0
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 0
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 0
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 0
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 0
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 0
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 0
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_405
timestamp 0
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 0
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 0
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 0
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 0
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 0
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 0
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 0
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 0
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 0
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 0
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 0
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 0
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 0
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 0
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 0
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 0
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 0
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 0
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 0
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 0
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 0
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 0
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 0
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 0
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 0
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 0
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_401
timestamp 0
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 0
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 0
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 0
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 0
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 0
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 0
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 0
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 0
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 0
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 0
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 0
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 0
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 0
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 0
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 0
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 0
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 0
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 0
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 0
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 0
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 0
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 0
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 0
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 0
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_405
timestamp 0
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 0
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 0
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 0
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 0
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 0
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 0
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 0
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 0
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 0
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 0
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 0
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 0
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 0
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 0
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 0
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 0
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 0
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 0
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 0
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 0
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 0
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 0
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 0
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 0
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 0
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 0
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_401
timestamp 0
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 0
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 0
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 0
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 0
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 0
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 0
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 0
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 0
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 0
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 0
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 0
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 0
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 0
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 0
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 0
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 0
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 0
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 0
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 0
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 0
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 0
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 0
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 0
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 0
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 0
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 0
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_405
timestamp 0
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 0
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 0
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 0
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 0
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 0
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 0
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 0
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 0
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 0
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 0
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 0
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 0
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 0
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 0
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 0
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 0
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 0
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 0
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 0
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 0
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 0
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 0
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 0
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 0
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 0
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 0
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_401
timestamp 0
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 0
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 0
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 0
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 0
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 0
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 0
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 0
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 0
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 0
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 0
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 0
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 0
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 0
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 0
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 0
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 0
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 0
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 0
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 0
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 0
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 0
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 0
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 0
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 0
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 0
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 0
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 0
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 0
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 0
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_405
timestamp 0
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 0
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 0
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 0
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 0
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 0
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 0
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 0
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 0
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 0
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 0
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 0
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 0
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 0
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 0
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 0
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 0
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 0
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 0
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 0
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 0
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 0
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 0
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 0
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 0
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 0
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 0
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_401
timestamp 0
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 0
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 0
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 0
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 0
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 0
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 0
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 0
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 0
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 0
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 0
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 0
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 0
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 0
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 0
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 0
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 0
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 0
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 0
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 0
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 0
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 0
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 0
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 0
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 0
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 0
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 0
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 0
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_405
timestamp 0
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 0
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 0
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 0
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 0
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 0
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 0
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 0
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 0
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 0
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 0
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 0
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 0
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 0
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 0
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 0
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 0
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 0
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 0
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 0
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 0
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 0
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 0
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 0
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 0
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_401
timestamp 0
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 0
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 0
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 0
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 0
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 0
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 0
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 0
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 0
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 0
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 0
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 0
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 0
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 0
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 0
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 0
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 0
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 0
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 0
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 0
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 0
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 0
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 0
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 0
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 0
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 0
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 0
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 0
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_405
timestamp 0
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 0
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 0
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 0
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 0
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 0
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 0
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 0
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 0
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 0
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 0
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 0
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 0
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 0
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 0
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 0
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 0
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 0
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 0
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 0
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 0
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 0
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 0
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 0
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 0
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 0
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_401
timestamp 0
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 0
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 0
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 0
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 0
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 0
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 0
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 0
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 0
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 0
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 0
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 0
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 0
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 0
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 0
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 0
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 0
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 0
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 0
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 0
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 0
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 0
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 0
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 0
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 0
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 0
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 0
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 0
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 0
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 0
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_405
timestamp 0
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 0
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 0
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 0
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 0
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 0
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 0
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 0
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 0
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 0
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 0
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 0
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 0
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 0
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 0
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 0
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 0
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 0
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 0
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 0
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 0
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 0
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 0
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 0
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 0
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 0
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 0
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 0
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 0
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_401
timestamp 0
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 0
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 0
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 0
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 0
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 0
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 0
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 0
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 0
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 0
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 0
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 0
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 0
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 0
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 0
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 0
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 0
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 0
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 0
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 0
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 0
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 0
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 0
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 0
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 0
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_361
timestamp 0
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 0
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 0
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 0
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 0
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_405
timestamp 0
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 0
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 0
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 0
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 0
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 0
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 0
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 0
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 0
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 0
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 0
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 0
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 0
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 0
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 0
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 0
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 0
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 0
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 0
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 0
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 0
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 0
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 0
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 0
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 0
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 0
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 0
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 0
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_401
timestamp 0
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 0
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 0
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 0
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 0
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 0
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 0
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 0
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 0
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 0
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 0
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 0
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 0
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 0
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 0
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 0
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 0
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 0
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 0
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 0
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 0
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 0
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_361
timestamp 0
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_373
timestamp 0
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_385
timestamp 0
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 0
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 0
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_405
timestamp 0
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 0
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 0
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 0
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 0
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 0
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 0
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 0
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 0
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 0
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 0
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 0
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 0
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 0
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 0
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 0
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 0
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 0
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 0
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 0
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 0
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 0
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 0
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 0
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 0
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 0
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 0
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 0
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 0
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_401
timestamp 0
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 0
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 0
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 0
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 0
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 0
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 0
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 0
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 0
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 0
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 0
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 0
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 0
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 0
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 0
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 0
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 0
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 0
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 0
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 0
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 0
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 0
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 0
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 0
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 0
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_361
timestamp 0
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 0
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_385
timestamp 0
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 0
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 0
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_405
timestamp 0
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 0
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 0
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 0
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 0
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 0
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 0
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 0
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 0
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 0
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 0
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 0
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 0
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 0
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 0
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 0
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 0
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 0
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 0
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 0
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 0
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 0
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 0
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 0
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 0
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 0
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 0
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 0
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 0
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 0
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 0
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_401
timestamp 0
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 0
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 0
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 0
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 0
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 0
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 0
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 0
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 0
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 0
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 0
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 0
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 0
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 0
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 0
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 0
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 0
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 0
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 0
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 0
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 0
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 0
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 0
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 0
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 0
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 0
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 0
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_361
timestamp 0
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_373
timestamp 0
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 0
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 0
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 0
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_405
timestamp 0
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 0
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 0
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 0
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 0
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 0
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 0
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 0
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 0
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 0
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 0
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 0
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 0
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 0
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 0
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 0
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 0
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 0
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 0
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 0
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 0
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 0
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 0
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 0
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 0
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 0
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 0
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 0
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 0
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 0
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 0
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 0
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 0
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 0
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 0
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_401
timestamp 0
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 0
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 0
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 0
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 0
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 0
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 0
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 0
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 0
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 0
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 0
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 0
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 0
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_193
timestamp 0
transform 1 0 18860 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_199
timestamp 0
transform 1 0 19412 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_209
timestamp 0
transform 1 0 20332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 0
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 0
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 0
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 0
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 0
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 0
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 0
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 0
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 0
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 0
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 0
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 0
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 0
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 0
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 0
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 0
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_385
timestamp 0
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 0
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 0
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_405
timestamp 0
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_7
timestamp 0
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_19
timestamp 0
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 0
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 0
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 0
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 0
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 0
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 0
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 0
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 0
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 0
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 0
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 0
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 0
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 0
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 0
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_197
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_218
timestamp 0
transform 1 0 21160 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_241
timestamp 0
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_249
timestamp 0
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 0
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 0
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 0
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 0
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 0
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 0
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 0
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 0
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 0
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 0
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 0
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 0
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 0
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 0
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 0
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_401
timestamp 0
transform 1 0 37996 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_6
timestamp 0
transform 1 0 1656 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_18
timestamp 0
transform 1 0 2760 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_30
timestamp 0
transform 1 0 3864 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_42
timestamp 0
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 0
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 0
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 0
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 0
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 0
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 0
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 0
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 0
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 0
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 0
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_181
timestamp 0
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_189
timestamp 0
transform 1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_220
timestamp 0
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 0
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 0
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 0
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 0
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 0
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 0
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 0
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 0
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 0
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 0
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 0
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 0
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 0
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 0
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 0
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 0
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 0
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 0
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_393
timestamp 0
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_401
timestamp 0
transform 1 0 37996 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_7
timestamp 0
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_19
timestamp 0
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 0
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 0
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 0
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 0
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 0
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 0
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 0
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 0
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 0
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 0
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_177
timestamp 0
transform 1 0 17388 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_185
timestamp 0
transform 1 0 18124 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_197
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_231
timestamp 0
transform 1 0 22356 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_243
timestamp 0
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 0
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 0
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 0
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 0
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 0
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 0
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 0
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 0
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 0
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 0
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 0
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 0
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 0
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 0
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 0
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 0
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_401
timestamp 0
transform 1 0 37996 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 0
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 0
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 0
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 0
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 0
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 0
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 0
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 0
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 0
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 0
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 0
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 0
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 0
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 0
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 0
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_193
timestamp 0
transform 1 0 18860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_216
timestamp 0
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 0
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 0
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 0
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 0
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 0
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 0
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 0
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 0
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 0
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 0
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 0
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 0
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 0
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 0
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 0
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 0
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 0
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 0
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_405
timestamp 0
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_6
timestamp 0
transform 1 0 1656 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_18
timestamp 0
transform 1 0 2760 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_26
timestamp 0
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 0
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 0
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 0
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 0
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 0
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 0
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 0
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 0
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 0
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 0
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 0
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 0
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 0
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 0
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 0
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 0
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 0
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 0
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 0
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 0
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 0
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 0
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 0
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 0
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 0
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 0
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 0
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 0
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 0
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 0
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 0
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 0
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 0
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_401
timestamp 0
transform 1 0 37996 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_7
timestamp 0
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_19
timestamp 0
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_31
timestamp 0
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_43
timestamp 0
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 0
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 0
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 0
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 0
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 0
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 0
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 0
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 0
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 0
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 0
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 0
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_181
timestamp 0
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_189
timestamp 0
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_211
timestamp 0
transform 1 0 20516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 0
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 0
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 0
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 0
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 0
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 0
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 0
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 0
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 0
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 0
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 0
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 0
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 0
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 0
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 0
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_373
timestamp 0
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 0
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 0
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_393
timestamp 0
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_401
timestamp 0
transform 1 0 37996 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 0
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 0
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 0
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 0
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 0
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 0
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 0
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 0
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 0
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 0
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 0
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 0
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 0
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 0
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 0
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 0
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 0
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 0
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 0
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 0
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 0
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 0
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 0
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 0
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 0
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 0
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 0
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 0
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 0
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 0
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 0
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 0
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 0
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 0
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 0
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 0
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 0
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_401
timestamp 0
transform 1 0 37996 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 0
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 0
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 0
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 0
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 0
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 0
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 0
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 0
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 0
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 0
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 0
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 0
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 0
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 0
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 0
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 0
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 0
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 0
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 0
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 0
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 0
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 0
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 0
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 0
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 0
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 0
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 0
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 0
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 0
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 0
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 0
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 0
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 0
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 0
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 0
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 0
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 0
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 0
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_405
timestamp 0
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 0
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 0
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 0
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 0
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 0
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 0
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 0
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 0
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 0
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 0
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 0
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 0
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 0
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 0
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 0
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 0
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 0
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 0
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 0
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 0
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 0
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 0
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 0
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 0
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 0
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 0
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 0
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 0
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 0
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 0
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 0
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 0
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 0
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 0
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 0
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 0
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_401
timestamp 0
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 0
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 0
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 0
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 0
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 0
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 0
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 0
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 0
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 0
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 0
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 0
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 0
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 0
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 0
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 0
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 0
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 0
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 0
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 0
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 0
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 0
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 0
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 0
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 0
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 0
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 0
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 0
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 0
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 0
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 0
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 0
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 0
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 0
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 0
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 0
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_361
timestamp 0
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_373
timestamp 0
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_385
timestamp 0
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 0
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 0
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_405
timestamp 0
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 0
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 0
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 0
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 0
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 0
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 0
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 0
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 0
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 0
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 0
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 0
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 0
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 0
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 0
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 0
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 0
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 0
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 0
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 0
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 0
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 0
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 0
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 0
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 0
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 0
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 0
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 0
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 0
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 0
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 0
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 0
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 0
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 0
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 0
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 0
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 0
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 0
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 0
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 0
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_401
timestamp 0
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 0
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 0
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 0
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 0
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 0
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 0
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 0
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 0
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 0
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 0
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 0
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 0
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 0
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 0
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 0
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 0
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 0
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 0
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 0
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 0
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 0
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 0
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 0
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 0
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 0
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 0
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 0
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 0
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 0
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 0
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 0
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 0
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 0
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 0
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 0
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 0
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 0
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 0
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 0
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 0
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_405
timestamp 0
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 0
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 0
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 0
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 0
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 0
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 0
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 0
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 0
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 0
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 0
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 0
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 0
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 0
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 0
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 0
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 0
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 0
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 0
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 0
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 0
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 0
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 0
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 0
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 0
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 0
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 0
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 0
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 0
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 0
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 0
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 0
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 0
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 0
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 0
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 0
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 0
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 0
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 0
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 0
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 0
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 0
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 0
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_401
timestamp 0
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 0
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 0
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 0
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 0
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 0
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 0
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 0
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 0
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 0
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 0
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 0
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 0
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 0
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 0
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 0
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 0
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 0
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 0
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 0
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 0
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 0
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 0
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 0
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 0
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 0
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 0
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 0
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 0
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 0
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 0
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 0
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 0
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 0
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 0
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 0
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 0
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 0
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 0
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 0
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 0
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 0
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 0
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 0
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_405
timestamp 0
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 0
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 0
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 0
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 0
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 0
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 0
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 0
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 0
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 0
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 0
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 0
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 0
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 0
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 0
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 0
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 0
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 0
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 0
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 0
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 0
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 0
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 0
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 0
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 0
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 0
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 0
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 0
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 0
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 0
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 0
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 0
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 0
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 0
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 0
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 0
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 0
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 0
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 0
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 0
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 0
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 0
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 0
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_401
timestamp 0
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 0
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 0
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 0
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 0
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 0
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 0
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 0
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 0
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 0
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 0
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 0
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 0
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 0
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 0
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 0
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 0
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 0
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 0
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 0
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 0
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 0
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 0
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 0
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 0
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 0
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 0
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 0
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 0
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 0
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 0
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 0
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 0
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 0
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 0
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 0
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 0
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 0
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 0
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 0
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 0
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 0
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 0
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 0
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_405
timestamp 0
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 0
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 0
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 0
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 0
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 0
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 0
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 0
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 0
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 0
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 0
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 0
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 0
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 0
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 0
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 0
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 0
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 0
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 0
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 0
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 0
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 0
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 0
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 0
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 0
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 0
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 0
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 0
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 0
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 0
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 0
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 0
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 0
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 0
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 0
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 0
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 0
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 0
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 0
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 0
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 0
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 0
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 0
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_401
timestamp 0
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 0
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 0
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 0
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 0
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 0
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 0
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 0
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 0
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 0
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 0
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 0
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 0
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 0
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 0
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 0
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 0
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 0
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 0
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 0
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 0
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 0
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 0
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 0
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 0
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 0
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 0
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 0
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 0
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 0
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 0
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 0
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 0
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 0
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 0
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 0
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 0
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 0
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 0
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 0
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 0
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 0
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 0
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 0
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_405
timestamp 0
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 0
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 0
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 0
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 0
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 0
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 0
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 0
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 0
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 0
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 0
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 0
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 0
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 0
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 0
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 0
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 0
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 0
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 0
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 0
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 0
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 0
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 0
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 0
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 0
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 0
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 0
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 0
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 0
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 0
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 0
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 0
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 0
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 0
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 0
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 0
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 0
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 0
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 0
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 0
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 0
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 0
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 0
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_401
timestamp 0
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 0
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 0
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 0
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 0
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 0
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 0
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 0
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 0
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 0
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 0
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 0
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 0
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 0
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 0
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 0
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 0
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 0
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 0
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 0
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 0
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 0
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 0
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 0
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 0
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 0
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 0
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 0
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 0
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 0
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 0
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 0
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 0
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 0
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 0
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 0
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 0
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 0
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 0
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 0
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 0
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 0
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 0
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 0
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_405
timestamp 0
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 0
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 0
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 0
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 0
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 0
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 0
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 0
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 0
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 0
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 0
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 0
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 0
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 0
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 0
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 0
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 0
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 0
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 0
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 0
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 0
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 0
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 0
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 0
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 0
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 0
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 0
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 0
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 0
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 0
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 0
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 0
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 0
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 0
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 0
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 0
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 0
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 0
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 0
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 0
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 0
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 0
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 0
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_401
timestamp 0
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 0
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 0
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 0
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 0
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 0
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 0
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 0
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 0
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 0
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 0
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 0
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 0
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 0
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 0
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 0
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 0
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 0
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 0
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 0
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 0
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 0
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 0
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 0
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 0
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 0
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 0
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 0
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 0
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 0
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 0
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 0
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 0
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 0
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 0
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 0
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 0
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 0
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 0
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 0
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 0
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 0
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 0
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 0
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_405
timestamp 0
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 0
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 0
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 0
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 0
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 0
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 0
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 0
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 0
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 0
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 0
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 0
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 0
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 0
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 0
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 0
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 0
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 0
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 0
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 0
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 0
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 0
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 0
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 0
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 0
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 0
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 0
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 0
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 0
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 0
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 0
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 0
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 0
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 0
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 0
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 0
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 0
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 0
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 0
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 0
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 0
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 0
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 0
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_401
timestamp 0
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 0
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 0
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 0
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 0
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 0
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 0
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 0
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 0
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 0
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 0
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 0
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 0
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 0
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 0
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 0
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 0
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 0
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 0
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 0
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 0
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 0
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 0
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 0
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 0
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 0
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 0
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 0
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 0
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 0
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 0
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 0
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 0
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 0
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 0
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 0
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 0
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 0
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 0
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 0
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 0
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 0
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 0
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 0
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_405
timestamp 0
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 0
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 0
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 0
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 0
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 0
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 0
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 0
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 0
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 0
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 0
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 0
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 0
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 0
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 0
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 0
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 0
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 0
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 0
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 0
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 0
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 0
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 0
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 0
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 0
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 0
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 0
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 0
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 0
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 0
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 0
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 0
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 0
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 0
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 0
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 0
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 0
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 0
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 0
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 0
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 0
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 0
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 0
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_401
timestamp 0
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 0
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 0
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 0
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 0
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 0
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 0
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 0
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 0
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 0
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 0
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 0
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 0
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 0
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 0
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 0
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 0
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 0
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 0
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 0
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 0
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 0
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 0
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 0
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 0
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 0
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 0
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 0
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 0
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 0
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 0
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 0
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 0
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 0
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 0
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 0
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 0
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 0
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 0
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 0
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 0
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 0
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 0
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 0
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_405
timestamp 0
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 0
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 0
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 0
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 0
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 0
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 0
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 0
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 0
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 0
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 0
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 0
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 0
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 0
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 0
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 0
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 0
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 0
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 0
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 0
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 0
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 0
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 0
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 0
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 0
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 0
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 0
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 0
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 0
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 0
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 0
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 0
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 0
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 0
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 0
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 0
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 0
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 0
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 0
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 0
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 0
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 0
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 0
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_401
timestamp 0
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 0
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 0
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 0
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 0
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 0
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 0
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 0
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 0
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 0
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 0
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 0
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 0
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 0
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 0
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 0
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 0
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 0
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 0
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 0
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 0
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 0
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 0
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 0
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 0
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 0
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 0
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 0
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 0
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 0
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 0
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 0
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 0
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 0
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 0
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 0
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 0
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 0
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 0
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 0
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 0
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 0
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 0
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 0
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_405
timestamp 0
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 0
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 0
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 0
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 0
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 0
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 0
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 0
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 0
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 0
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 0
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 0
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 0
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 0
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 0
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 0
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 0
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 0
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 0
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 0
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 0
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 0
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 0
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 0
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 0
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 0
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 0
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 0
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 0
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 0
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 0
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 0
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 0
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 0
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 0
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 0
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 0
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 0
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 0
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 0
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 0
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 0
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 0
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_401
timestamp 0
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 0
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 0
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 0
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 0
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 0
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 0
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 0
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 0
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 0
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 0
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 0
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 0
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 0
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 0
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 0
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 0
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 0
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 0
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 0
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 0
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 0
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 0
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 0
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 0
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 0
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 0
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 0
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 0
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 0
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 0
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 0
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 0
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 0
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 0
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 0
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 0
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 0
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 0
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 0
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 0
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 0
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 0
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 0
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_405
timestamp 0
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 0
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 0
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 0
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 0
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 0
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 0
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 0
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 0
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 0
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 0
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 0
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 0
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 0
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 0
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 0
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 0
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 0
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 0
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 0
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 0
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 0
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 0
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 0
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 0
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 0
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 0
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 0
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 0
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 0
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 0
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 0
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 0
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 0
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 0
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 0
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 0
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 0
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 0
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 0
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 0
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 0
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 0
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_401
timestamp 0
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 0
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 0
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 0
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 0
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 0
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 0
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 0
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 0
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 0
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 0
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 0
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 0
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 0
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 0
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 0
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 0
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 0
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 0
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 0
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 0
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 0
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 0
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 0
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 0
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 0
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 0
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 0
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 0
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 0
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 0
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 0
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 0
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 0
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 0
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 0
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 0
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 0
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 0
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 0
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 0
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 0
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 0
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 0
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_405
timestamp 0
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 0
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 0
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 0
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 0
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 0
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 0
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 0
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 0
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 0
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 0
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 0
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 0
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 0
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 0
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 0
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 0
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 0
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 0
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 0
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 0
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 0
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 0
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 0
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 0
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 0
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 0
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 0
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 0
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 0
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 0
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 0
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 0
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 0
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 0
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 0
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 0
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 0
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 0
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 0
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 0
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 0
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 0
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_401
timestamp 0
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 0
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 0
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 0
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 0
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 0
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 0
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 0
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 0
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 0
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 0
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 0
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 0
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 0
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 0
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 0
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 0
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 0
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 0
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 0
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 0
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 0
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 0
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 0
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 0
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 0
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 0
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 0
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 0
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 0
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 0
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 0
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 0
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 0
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 0
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 0
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 0
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 0
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 0
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 0
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 0
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 0
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 0
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 0
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_405
timestamp 0
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 0
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 0
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 0
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 0
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 0
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_53
timestamp 0
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_57
timestamp 0
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_69
timestamp 0
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_81
timestamp 0
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 0
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 0
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_109
timestamp 0
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_113
timestamp 0
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 0
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 0
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 0
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 0
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_165
timestamp 0
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_169
timestamp 0
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_181
timestamp 0
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 0
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 0
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 0
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_221
timestamp 0
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_225
timestamp 0
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_237
timestamp 0
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_249
timestamp 0
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 0
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 0
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_277
timestamp 0
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_281
timestamp 0
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_293
timestamp 0
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_305
timestamp 0
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 0
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 0
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_333
timestamp 0
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_337
timestamp 0
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_349
timestamp 0
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_361
timestamp 0
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 0
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 0
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_389
timestamp 0
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_393
timestamp 0
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_405
timestamp 0
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  out_sky130_fd_sc_hd__buf_1_X_1
timestamp 0
transform 1 0 20700 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  out_sky130_fd_sc_hd__buf_1_X_2
timestamp 0
transform 1 0 21804 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  out_sky130_fd_sc_hd__buf_1_X_3
timestamp 0
transform 1 0 18768 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  out_sky130_fd_sc_hd__buf_1_X_4
timestamp 0
transform 1 0 20424 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  out_sky130_fd_sc_hd__buf_1_X_5
timestamp 0
transform -1 0 19504 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  out_sky130_fd_sc_hd__buf_1_X
timestamp 0
transform 1 0 22080 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  out_sky130_fd_sc_hd__buf_1_X_6
timestamp 0
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_2  out_sky130_fd_sc_hd__nor4b_2_Y
timestamp 0
transform -1 0 20424 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  output4
timestamp 0
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output5
timestamp 0
transform 1 0 38272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output6
timestamp 0
transform -1 0 1656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output7
timestamp 0
transform 1 0 38272 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output8
timestamp 0
transform 1 0 38272 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output9
timestamp 0
transform 1 0 38272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output10
timestamp 0
transform 1 0 38272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output11
timestamp 0
transform 1 0 38272 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_65
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_66
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_67
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_68
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_69
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_70
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_71
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_72
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_73
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_74
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_75
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_76
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_77
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_78
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_79
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_80
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_81
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_82
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_83
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_84
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_85
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_86
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_87
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_88
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_89
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_90
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_91
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_92
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_93
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 0
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_94
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 0
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_95
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 0
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_96
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 0
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_97
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 0
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_98
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 0
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_99
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 0
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_100
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 0
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_101
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 0
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_102
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 0
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_103
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 0
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_104
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 0
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_105
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 0
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_106
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 0
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_107
timestamp 0
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 0
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_108
timestamp 0
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 0
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_109
timestamp 0
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 0
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_110
timestamp 0
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 0
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_111
timestamp 0
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 0
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_112
timestamp 0
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 0
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_113
timestamp 0
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 0
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_114
timestamp 0
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 0
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_115
timestamp 0
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 0
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_116
timestamp 0
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 0
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_117
timestamp 0
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 0
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_118
timestamp 0
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 0
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_119
timestamp 0
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 0
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_120
timestamp 0
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 0
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_121
timestamp 0
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 0
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_122
timestamp 0
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 0
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_123
timestamp 0
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 0
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_124
timestamp 0
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 0
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_125
timestamp 0
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 0
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_126
timestamp 0
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 0
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_127
timestamp 0
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 0
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_128
timestamp 0
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 0
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_129
timestamp 0
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 0
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 0
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 0
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 0
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 0
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 0
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_143
timestamp 0
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_144
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_145
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_146
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_147
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_148
timestamp 0
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_149
timestamp 0
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_150
timestamp 0
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_151
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_152
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_153
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_154
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_155
timestamp 0
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_156
timestamp 0
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_157
timestamp 0
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_158
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_159
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_160
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_161
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_162
timestamp 0
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_163
timestamp 0
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_164
timestamp 0
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_165
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_166
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_167
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_168
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_169
timestamp 0
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_170
timestamp 0
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_171
timestamp 0
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_172
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_173
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_174
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_175
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_176
timestamp 0
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_177
timestamp 0
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_178
timestamp 0
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_179
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_180
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_181
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_182
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_183
timestamp 0
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_184
timestamp 0
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_185
timestamp 0
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_186
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_187
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_188
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_189
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_190
timestamp 0
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_191
timestamp 0
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_192
timestamp 0
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_193
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_194
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_195
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_196
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_197
timestamp 0
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_198
timestamp 0
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_199
timestamp 0
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_200
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_201
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_202
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_203
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_204
timestamp 0
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_205
timestamp 0
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_206
timestamp 0
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_207
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_208
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_209
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_210
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_211
timestamp 0
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_212
timestamp 0
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_213
timestamp 0
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_214
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_215
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_216
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_217
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_218
timestamp 0
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_219
timestamp 0
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_220
timestamp 0
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_221
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_222
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_223
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_224
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_225
timestamp 0
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_226
timestamp 0
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_227
timestamp 0
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_228
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_229
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_230
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_231
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_232
timestamp 0
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_233
timestamp 0
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_234
timestamp 0
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_235
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_236
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_237
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_238
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_239
timestamp 0
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_240
timestamp 0
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_241
timestamp 0
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_242
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_243
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_244
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_245
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_246
timestamp 0
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_247
timestamp 0
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_248
timestamp 0
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_249
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_250
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_251
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_252
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_253
timestamp 0
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_254
timestamp 0
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_255
timestamp 0
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_256
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_257
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_258
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_259
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_260
timestamp 0
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_261
timestamp 0
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_262
timestamp 0
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_263
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_264
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_265
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_266
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_267
timestamp 0
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_268
timestamp 0
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_269
timestamp 0
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_270
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_271
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_272
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_273
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_274
timestamp 0
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_275
timestamp 0
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_276
timestamp 0
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_277
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_278
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_279
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_280
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_281
timestamp 0
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_282
timestamp 0
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_283
timestamp 0
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_284
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_285
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_286
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_287
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_288
timestamp 0
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_289
timestamp 0
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_290
timestamp 0
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_291
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_292
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_293
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_294
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_295
timestamp 0
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_296
timestamp 0
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_297
timestamp 0
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_298
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_299
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_300
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_301
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_302
timestamp 0
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_303
timestamp 0
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_304
timestamp 0
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_305
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_306
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_307
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_308
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_309
timestamp 0
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_310
timestamp 0
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_311
timestamp 0
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_312
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_313
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_314
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_315
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_316
timestamp 0
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_317
timestamp 0
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_318
timestamp 0
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_319
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_320
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_321
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_322
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_323
timestamp 0
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_324
timestamp 0
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_325
timestamp 0
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_326
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_327
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_328
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_329
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_330
timestamp 0
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_331
timestamp 0
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_332
timestamp 0
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_333
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_334
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_335
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_336
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_337
timestamp 0
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_338
timestamp 0
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_339
timestamp 0
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_340
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_341
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_342
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_343
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_344
timestamp 0
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_345
timestamp 0
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_346
timestamp 0
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_347
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_348
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_349
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_350
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_351
timestamp 0
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_352
timestamp 0
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_353
timestamp 0
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_354
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_355
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_356
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_357
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_358
timestamp 0
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_359
timestamp 0
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_360
timestamp 0
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_361
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_362
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_363
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_364
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_365
timestamp 0
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_366
timestamp 0
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_367
timestamp 0
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_368
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_369
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_370
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_371
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_372
timestamp 0
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_373
timestamp 0
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_374
timestamp 0
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_375
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_376
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_377
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_378
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_379
timestamp 0
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_380
timestamp 0
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_381
timestamp 0
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_382
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_383
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_384
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_385
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_386
timestamp 0
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_387
timestamp 0
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_388
timestamp 0
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_389
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_390
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_391
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_392
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_393
timestamp 0
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_394
timestamp 0
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_395
timestamp 0
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_396
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_397
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_398
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_399
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_400
timestamp 0
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_401
timestamp 0
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_402
timestamp 0
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_403
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_404
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_405
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_406
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_407
timestamp 0
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_408
timestamp 0
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_409
timestamp 0
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_410
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_411
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_412
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_413
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_414
timestamp 0
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_415
timestamp 0
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_416
timestamp 0
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_417
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_418
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_419
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_420
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_421
timestamp 0
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_422
timestamp 0
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_423
timestamp 0
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_424
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_425
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_426
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_427
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_428
timestamp 0
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_429
timestamp 0
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_430
timestamp 0
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_431
timestamp 0
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_432
timestamp 0
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_433
timestamp 0
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_434
timestamp 0
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_435
timestamp 0
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_436
timestamp 0
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_437
timestamp 0
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_438
timestamp 0
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_439
timestamp 0
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_440
timestamp 0
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_441
timestamp 0
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_442
timestamp 0
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_443
timestamp 0
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_444
timestamp 0
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_445
timestamp 0
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_446
timestamp 0
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_447
timestamp 0
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_448
timestamp 0
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_449
timestamp 0
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_450
timestamp 0
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_451
timestamp 0
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_452
timestamp 0
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_453
timestamp 0
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_454
timestamp 0
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_455
timestamp 0
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_456
timestamp 0
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_457
timestamp 0
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_458
timestamp 0
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_459
timestamp 0
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_460
timestamp 0
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_461
timestamp 0
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_462
timestamp 0
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_463
timestamp 0
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_464
timestamp 0
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_465
timestamp 0
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_466
timestamp 0
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_467
timestamp 0
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_468
timestamp 0
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_469
timestamp 0
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_470
timestamp 0
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_471
timestamp 0
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_472
timestamp 0
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_473
timestamp 0
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_474
timestamp 0
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_475
timestamp 0
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_476
timestamp 0
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_477
timestamp 0
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_478
timestamp 0
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_479
timestamp 0
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_480
timestamp 0
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_481
timestamp 0
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_482
timestamp 0
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_483
timestamp 0
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_484
timestamp 0
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_485
timestamp 0
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_486
timestamp 0
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_487
timestamp 0
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_488
timestamp 0
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_489
timestamp 0
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_490
timestamp 0
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_491
timestamp 0
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_492
timestamp 0
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_493
timestamp 0
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_494
timestamp 0
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_495
timestamp 0
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_496
timestamp 0
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_497
timestamp 0
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_498
timestamp 0
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_499
timestamp 0
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_500
timestamp 0
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_501
timestamp 0
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_502
timestamp 0
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_503
timestamp 0
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_504
timestamp 0
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_505
timestamp 0
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_506
timestamp 0
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_507
timestamp 0
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_508
timestamp 0
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_509
timestamp 0
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_510
timestamp 0
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_511
timestamp 0
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_512
timestamp 0
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_513
timestamp 0
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_514
timestamp 0
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_515
timestamp 0
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_516
timestamp 0
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_517
timestamp 0
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_518
timestamp 0
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_519
timestamp 0
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_520
timestamp 0
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_521
timestamp 0
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_522
timestamp 0
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_523
timestamp 0
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_524
timestamp 0
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_525
timestamp 0
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_526
timestamp 0
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_527
timestamp 0
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_528
timestamp 0
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_529
timestamp 0
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_530
timestamp 0
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_531
timestamp 0
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_532
timestamp 0
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_533
timestamp 0
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_534
timestamp 0
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_535
timestamp 0
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_536
timestamp 0
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_537
timestamp 0
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_538
timestamp 0
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_539
timestamp 0
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_540
timestamp 0
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_541
timestamp 0
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_542
timestamp 0
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_543
timestamp 0
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_544
timestamp 0
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_545
timestamp 0
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_546
timestamp 0
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_547
timestamp 0
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_548
timestamp 0
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_549
timestamp 0
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_550
timestamp 0
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_551
timestamp 0
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_552
timestamp 0
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_553
timestamp 0
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_554
timestamp 0
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_555
timestamp 0
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_556
timestamp 0
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_557
timestamp 0
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_558
timestamp 0
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_559
timestamp 0
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_560
timestamp 0
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_561
timestamp 0
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_562
timestamp 0
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_563
timestamp 0
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_564
timestamp 0
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_565
timestamp 0
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_566
timestamp 0
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_567
timestamp 0
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_568
timestamp 0
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_569
timestamp 0
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_570
timestamp 0
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_571
timestamp 0
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_572
timestamp 0
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_573
timestamp 0
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_574
timestamp 0
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_575
timestamp 0
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_576
timestamp 0
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_577
timestamp 0
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_578
timestamp 0
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_579
timestamp 0
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_580
timestamp 0
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_581
timestamp 0
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_582
timestamp 0
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_583
timestamp 0
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_584
timestamp 0
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_585
timestamp 0
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_586
timestamp 0
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_587
timestamp 0
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_588
timestamp 0
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_589
timestamp 0
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_590
timestamp 0
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_591
timestamp 0
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_592
timestamp 0
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_593
timestamp 0
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_594
timestamp 0
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_595
timestamp 0
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_596
timestamp 0
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_597
timestamp 0
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_598
timestamp 0
transform 1 0 37168 0 1 36992
box -38 -48 130 592
<< labels >>
rlabel metal1 s 19964 36992 19964 36992 4 VGND
rlabel metal1 s 19964 37536 19964 37536 4 VPWR
rlabel metal2 s 21758 19618 21758 19618 4 clk
rlabel metal1 s 20470 20468 20470 20468 4 clk_sky130_fd_sc_hd__and4b_2_B_X
rlabel metal1 s 20470 19822 20470 19822 4 clk_sky130_fd_sc_hd__and4b_2_C_X
rlabel metal1 s 20470 18394 20470 18394 4 clk_sky130_fd_sc_hd__and4b_2_D_X
rlabel metal2 s 20470 19244 20470 19244 4 clknet_0_clk
rlabel metal2 s 19826 21148 19826 21148 4 clknet_1_0__leaf_clk
rlabel metal1 s 21804 18598 21804 18598 4 clknet_1_1__leaf_clk
rlabel metal3 s 820 21148 820 21148 4 in[0]
rlabel metal3 s 820 19788 820 19788 4 in[1]
rlabel metal3 s 820 18428 820 18428 4 in[2]
rlabel metal2 s 1610 21216 1610 21216 4 net1
rlabel metal2 s 38318 20910 38318 20910 4 net10
rlabel metal2 s 34546 20434 34546 20434 4 net11
rlabel metal2 s 19550 20162 19550 20162 4 net2
rlabel metal2 s 18630 19278 18630 19278 4 net3
rlabel metal1 s 19642 19380 19642 19380 4 net4
rlabel metal1 s 21666 19448 21666 19448 4 net5
rlabel metal2 s 15226 20740 15226 20740 4 net6
rlabel metal1 s 20654 20264 20654 20264 4 net7
rlabel metal2 s 18998 19431 18998 19431 4 net8
rlabel metal1 s 22034 19720 22034 19720 4 net9
rlabel metal3 s 1050 19108 1050 19108 4 out[0]
rlabel metal1 s 38686 20026 38686 20026 4 out[1]
rlabel metal3 s 0 20408 800 20528 4 out[2]
port 9 nsew
rlabel metal3 s 38502 21845 38502 21845 4 out[3]
rlabel metal3 s 38502 19125 38502 19125 4 out[4]
rlabel metal2 s 38502 18513 38502 18513 4 out[5]
rlabel metal2 s 38502 21233 38502 21233 4 out[6]
rlabel metal1 s 38778 20774 38778 20774 4 out[7]
rlabel metal1 s 18906 19346 18906 19346 4 out_sky130_fd_sc_hd__buf_1_X_3_A
rlabel metal1 s 19596 18802 19596 18802 4 out_sky130_fd_sc_hd__buf_1_X_5_A
rlabel metal1 s 19228 19346 19228 19346 4 out_sky130_fd_sc_hd__buf_1_X_6_A
rlabel metal1 s 21666 18938 21666 18938 4 out_sky130_fd_sc_hd__buf_1_X_A
flabel metal5 s 1056 33676 38872 33996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 28676 38872 28996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 23676 38872 23996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 18676 38872 18996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 13676 38872 13996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8676 38872 8996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3676 38872 3996 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 37604 2128 37924 37584 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 32604 2128 32924 37584 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 27604 2128 27924 37584 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 22604 2128 22924 37584 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 17604 2128 17924 37584 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 12604 2128 12924 37584 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7604 2128 7924 37584 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2604 2128 2924 37584 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 33016 38872 33336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 28016 38872 28336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 23016 38872 23336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 18016 38872 18336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 13016 38872 13336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 8016 38872 8336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3016 38872 3336 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 36944 2128 37264 37584 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 31944 2128 32264 37584 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 26944 2128 27264 37584 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 21944 2128 22264 37584 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 16944 2128 17264 37584 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 11944 2128 12264 37584 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 6944 2128 7264 37584 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1944 2128 2264 37584 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 39200 17688 40000 17808 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 0 21088 800 21208 0 FreeSans 600 0 0 0 in[0]
port 4 nsew
flabel metal3 s 0 19728 800 19848 0 FreeSans 600 0 0 0 in[1]
port 5 nsew
flabel metal3 s 0 18368 800 18488 0 FreeSans 600 0 0 0 in[2]
port 6 nsew
flabel metal3 s 0 19048 800 19168 0 FreeSans 600 0 0 0 out[0]
port 7 nsew
flabel metal3 s 39200 19728 40000 19848 0 FreeSans 600 0 0 0 out[1]
port 8 nsew
flabel metal3 s 400 20468 400 20468 0 FreeSans 600 0 0 0 out[2]
flabel metal3 s 39200 21768 40000 21888 0 FreeSans 600 0 0 0 out[3]
port 10 nsew
flabel metal3 s 39200 19048 40000 19168 0 FreeSans 600 0 0 0 out[4]
port 11 nsew
flabel metal3 s 39200 18368 40000 18488 0 FreeSans 600 0 0 0 out[5]
port 12 nsew
flabel metal3 s 39200 21088 40000 21208 0 FreeSans 600 0 0 0 out[6]
port 13 nsew
flabel metal3 s 39200 20408 40000 20528 0 FreeSans 600 0 0 0 out[7]
port 14 nsew
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
