magic
tech sky130A
magscale 1 2
timestamp 1698989880
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 934 2128 39086 37584
<< obsm2 >>
rect 938 2139 39082 37573
<< metal3 >>
rect 39200 21768 40000 21888
rect 0 21088 800 21208
rect 39200 21088 40000 21208
rect 0 20408 800 20528
rect 39200 20408 40000 20528
rect 0 19728 800 19848
rect 39200 19728 40000 19848
rect 0 19048 800 19168
rect 39200 19048 40000 19168
rect 0 18368 800 18488
rect 39200 18368 40000 18488
rect 39200 17688 40000 17808
<< obsm3 >>
rect 798 21968 39200 37569
rect 798 21688 39120 21968
rect 798 21288 39200 21688
rect 880 21008 39120 21288
rect 798 20608 39200 21008
rect 880 20328 39120 20608
rect 798 19928 39200 20328
rect 880 19648 39120 19928
rect 798 19248 39200 19648
rect 880 18968 39120 19248
rect 798 18568 39200 18968
rect 880 18288 39120 18568
rect 798 17888 39200 18288
rect 798 17608 39120 17888
rect 798 2143 39200 17608
<< metal4 >>
rect 1944 2128 2264 37584
rect 2604 2128 2924 37584
rect 6944 2128 7264 37584
rect 7604 2128 7924 37584
rect 11944 2128 12264 37584
rect 12604 2128 12924 37584
rect 16944 2128 17264 37584
rect 17604 2128 17924 37584
rect 21944 2128 22264 37584
rect 22604 2128 22924 37584
rect 26944 2128 27264 37584
rect 27604 2128 27924 37584
rect 31944 2128 32264 37584
rect 32604 2128 32924 37584
rect 36944 2128 37264 37584
rect 37604 2128 37924 37584
<< metal5 >>
rect 1056 33676 38872 33996
rect 1056 33016 38872 33336
rect 1056 28676 38872 28996
rect 1056 28016 38872 28336
rect 1056 23676 38872 23996
rect 1056 23016 38872 23336
rect 1056 18676 38872 18996
rect 1056 18016 38872 18336
rect 1056 13676 38872 13996
rect 1056 13016 38872 13336
rect 1056 8676 38872 8996
rect 1056 8016 38872 8336
rect 1056 3676 38872 3996
rect 1056 3016 38872 3336
<< labels >>
rlabel metal4 s 2604 2128 2924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7604 2128 7924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12604 2128 12924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17604 2128 17924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 22604 2128 22924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27604 2128 27924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 32604 2128 32924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37604 2128 37924 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3676 38872 3996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8676 38872 8996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 13676 38872 13996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 18676 38872 18996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 23676 38872 23996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 28676 38872 28996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 33676 38872 33996 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6944 2128 7264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11944 2128 12264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16944 2128 17264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 21944 2128 22264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 26944 2128 27264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 31944 2128 32264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 36944 2128 37264 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3016 38872 3336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8016 38872 8336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 13016 38872 13336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 18016 38872 18336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 23016 38872 23336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 28016 38872 28336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 33016 38872 33336 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 39200 17688 40000 17808 6 clk
port 3 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 in[0]
port 4 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 in[1]
port 5 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 in[2]
port 6 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 out[0]
port 7 nsew signal output
rlabel metal3 s 39200 19728 40000 19848 6 out[1]
port 8 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 out[2]
port 9 nsew signal output
rlabel metal3 s 39200 21768 40000 21888 6 out[3]
port 10 nsew signal output
rlabel metal3 s 39200 19048 40000 19168 6 out[4]
port 11 nsew signal output
rlabel metal3 s 39200 18368 40000 18488 6 out[5]
port 12 nsew signal output
rlabel metal3 s 39200 21088 40000 21208 6 out[6]
port 13 nsew signal output
rlabel metal3 s 39200 20408 40000 20528 6 out[7]
port 14 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 938330
string GDS_FILE /openlane/openlane/pes_decoder/runs/RUN_CHECK/results/signoff/pes_decoder.magic.gds
string GDS_START 74440
<< end >>

